* NGSPICE file created from SPM_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

.subckt SPM_example VGND VPWR io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2106_ clknet_leaf_11_wb_clk_i _0393_ _0206_ VGND VGND VPWR VPWR Y\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2037_ clknet_leaf_5_wb_clk_i _0324_ _0170_ VGND VGND VPWR VPWR P0\[58\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1270_ CNT\[1\] CNT\[0\] CNT\[2\] VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__and3_1
XFILLER_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0985_ net49 Y\[22\] _0799_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__mux2_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1606_ _0594_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__inv_2
X_1537_ _0587_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1468_ _0570_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__nor2_1
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_260 VGND VGND VPWR VPWR SPM_example_260/HI la_data_out[74] sky130_fd_sc_hd__conb_1
XFILLER_67_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1399_ spm.csa0.sc spm.csa0.y VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__nor2_1
XSPM_example_271 VGND VGND VPWR VPWR SPM_example_271/HI la_data_out[85] sky130_fd_sc_hd__conb_1
XFILLER_110_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_282 VGND VGND VPWR VPWR SPM_example_282/HI la_data_out[96] sky130_fd_sc_hd__conb_1
XFILLER_132_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_293 VGND VGND VPWR VPWR SPM_example_293/HI la_data_out[107] sky130_fd_sc_hd__conb_1
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1322_ _0472_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nor2_1
XFILLER_96_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1253_ net61 spm.x\[4\] _0421_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1184_ _0925_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0968_ _0785_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__buf_4
XFILLER_118_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ clknet_leaf_20_wb_clk_i _0236_ _0073_ VGND VGND VPWR VPWR spm.x\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1871_ _0761_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__inv_2
XFILLER_187_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1305_ _0453_ spm.x\[15\] VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__nand2_1
XFILLER_57_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1236_ net38 spm.x\[12\] _0410_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1167_ P0\[11\] P0\[12\] _0914_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__mux2_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1098_ _0880_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2070_ clknet_leaf_6_wb_clk_i _0357_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_2
XFILLER_94_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1021_ _0834_ Y\[12\] _0817_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__mux2_1
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ clknet_leaf_18_wb_clk_i _0027_ _0056_ VGND VGND VPWR VPWR spm.genblk1\[6\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1854_ _0759_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__inv_2
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1785_ Y\[22\] _0700_ _0682_ _0716_ _0692_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__a221o_1
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2337_ net139 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_111_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1219_ _0411_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clknet_2_3__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_5 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1570_ _0590_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
XFILLER_67_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2122_ clknet_leaf_12_wb_clk_i spm.genblk1\[23\].csa.hsum2 _0222_ VGND VGND VPWR
+ VPWR spm.genblk1\[22\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2053_ clknet_leaf_23_wb_clk_i _0340_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_2
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1004_ _0823_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1906_ clknet_leaf_23_wb_clk_i spm.genblk1\[14\].csa.hsum2 _0039_ VGND VGND VPWR
+ VPWR spm.genblk1\[13\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_202_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1837_ _0598_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__inv_2
XFILLER_117_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1768_ P0\[51\] _0661_ _0662_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__o21a_1
XFILLER_117_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1699_ Y\[7\] _0779_ _0635_ _0644_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__a221o_1
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput75 net75 VGND VGND VPWR VPWR io_oeb[15] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VGND VGND VPWR VPWR io_oeb[25] sky130_fd_sc_hd__buf_2
Xoutput97 net97 VGND VGND VPWR VPWR io_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ _0596_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
XFILLER_132_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1553_ _0589_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
XFILLER_125_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1484_ net142 VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__clkbuf_4
XFILLER_141_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2105_ clknet_leaf_11_wb_clk_i _0392_ _0205_ VGND VGND VPWR VPWR Y\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2036_ clknet_leaf_4_wb_clk_i _0323_ _0169_ VGND VGND VPWR VPWR P0\[57\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_922 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0984_ _0809_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1605_ _0594_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__inv_2
XFILLER_133_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1536_ _0587_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_2
XFILLER_141_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout139 net140 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1467_ spm.genblk1\[20\].csa.sc spm.genblk1\[20\].csa.y VGND VGND VPWR VPWR _0571_
+ sky130_fd_sc_hd__and2_1
XSPM_example_250 VGND VGND VPWR VPWR SPM_example_250/HI la_data_out[64] sky130_fd_sc_hd__conb_1
XFILLER_80_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1398_ _0524_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
XSPM_example_261 VGND VGND VPWR VPWR SPM_example_261/HI la_data_out[75] sky130_fd_sc_hd__conb_1
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_272 VGND VGND VPWR VPWR SPM_example_272/HI la_data_out[86] sky130_fd_sc_hd__conb_1
XSPM_example_283 VGND VGND VPWR VPWR SPM_example_283/HI la_data_out[97] sky130_fd_sc_hd__conb_1
XFILLER_110_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_294 VGND VGND VPWR VPWR SPM_example_294/HI la_data_out[108] sky130_fd_sc_hd__conb_1
XFILLER_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2019_ clknet_leaf_24_wb_clk_i _0306_ _0152_ VGND VGND VPWR VPWR P0\[40\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1321_ spm.genblk1\[12\].csa.sc spm.genblk1\[12\].csa.y VGND VGND VPWR VPWR _0473_
+ sky130_fd_sc_hd__and2_1
XFILLER_2_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1252_ _0428_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1183_ P0\[3\] P0\[4\] _0793_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__mux2_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0967_ _0797_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1519_ _0586_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__inv_2
XFILLER_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1870_ _0761_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__inv_2
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1304_ _0460_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nor2_1
XFILLER_96_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1235_ _0419_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1166_ _0916_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1097_ P0\[44\] P0\[45\] _0870_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__mux2_1
XFILLER_197_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1999_ clknet_leaf_3_wb_clk_i _0286_ _0132_ VGND VGND VPWR VPWR P0\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_140_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1020_ net37 Y\[11\] _0821_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__mux2_1
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ clknet_leaf_18_wb_clk_i spm.genblk1\[6\].csa.hsum2 _0055_ VGND VGND VPWR VPWR
+ spm.genblk1\[5\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1853_ _0759_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__inv_2
XFILLER_147_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1784_ spm.x\[22\] P0\[22\] _0397_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__mux2_1
XFILLER_116_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2336_ net139 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1218_ net48 spm.x\[21\] _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1149_ _0907_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2121_ clknet_leaf_8_wb_clk_i _0016_ _0221_ VGND VGND VPWR VPWR spm.genblk1\[24\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2052_ clknet_leaf_23_wb_clk_i _0339_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_2
XFILLER_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1003_ _0822_ Y\[18\] _0817_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__mux2_1
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1905_ clknet_leaf_1_wb_clk_i _0006_ _0038_ VGND VGND VPWR VPWR spm.genblk1\[15\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1836_ _0756_ _0757_ _0758_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a21o_1
XFILLER_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1767_ Y\[19\] _0700_ _0682_ _0701_ _0692_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a221o_1
XFILLER_190_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1698_ _0605_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__clkbuf_4
XFILLER_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2319_ net142 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput76 net76 VGND VGND VPWR VPWR io_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_122_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput87 net87 VGND VGND VPWR VPWR io_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_1_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput98 net98 VGND VGND VPWR VPWR io_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1621_ _0596_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__inv_2
XFILLER_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1552_ _0589_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
XFILLER_67_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1483_ _0453_ spm.x\[18\] _0580_ _0579_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a31o_1
XFILLER_119_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2104_ clknet_leaf_8_wb_clk_i _0391_ _0204_ VGND VGND VPWR VPWR Y\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2035_ clknet_leaf_4_wb_clk_i _0322_ _0168_ VGND VGND VPWR VPWR P0\[56\] sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1819_ _0742_ _0743_ _0744_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a21o_1
XFILLER_117_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0983_ _0808_ Y\[24\] _0794_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__mux2_1
XFILLER_186_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1604_ _0594_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__inv_2
X_1535_ _0587_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_2
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1466_ spm.genblk1\[20\].csa.sc spm.genblk1\[20\].csa.y VGND VGND VPWR VPWR _0570_
+ sky130_fd_sc_hd__nor2_1
XFILLER_141_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1397_ _0032_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__and2_1
XSPM_example_240 VGND VGND VPWR VPWR SPM_example_240/HI la_data_out[54] sky130_fd_sc_hd__conb_1
XSPM_example_251 VGND VGND VPWR VPWR SPM_example_251/HI la_data_out[65] sky130_fd_sc_hd__conb_1
XFILLER_110_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_262 VGND VGND VPWR VPWR SPM_example_262/HI la_data_out[76] sky130_fd_sc_hd__conb_1
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_273 VGND VGND VPWR VPWR SPM_example_273/HI la_data_out[87] sky130_fd_sc_hd__conb_1
XSPM_example_284 VGND VGND VPWR VPWR SPM_example_284/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_295 VGND VGND VPWR VPWR SPM_example_295/HI la_data_out[109] sky130_fd_sc_hd__conb_1
XFILLER_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2018_ clknet_leaf_24_wb_clk_i _0305_ _0151_ VGND VGND VPWR VPWR P0\[39\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1320_ spm.genblk1\[12\].csa.sc spm.genblk1\[12\].csa.y VGND VGND VPWR VPWR _0472_
+ sky130_fd_sc_hd__nor2_1
XFILLER_116_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1251_ net62 spm.x\[5\] _0421_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux2_1
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1182_ _0924_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_0966_ _0796_ Y\[29\] _0794_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__mux2_1
XFILLER_203_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1518_ _0582_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__buf_4
XFILLER_88_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1449_ spm.genblk1\[23\].csa.sc spm.genblk1\[23\].csa.y VGND VGND VPWR VPWR _0559_
+ sky130_fd_sc_hd__and2_1
XFILLER_96_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1303_ spm.genblk1\[15\].csa.sc spm.genblk1\[15\].csa.y VGND VGND VPWR VPWR _0461_
+ sky130_fd_sc_hd__and2_1
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1234_ net39 spm.x\[13\] _0410_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
XFILLER_49_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1165_ P0\[12\] P0\[13\] _0914_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__mux2_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1096_ _0879_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1998_ clknet_leaf_3_wb_clk_i _0285_ _0131_ VGND VGND VPWR VPWR P0\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_165_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0949_ net19 net20 net26 net22 VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__or4b_1
XFILLER_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1921_ clknet_leaf_18_wb_clk_i _0028_ _0054_ VGND VGND VPWR VPWR spm.genblk1\[7\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_203_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1852_ _0759_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__inv_2
XFILLER_124_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1783_ _0713_ _0714_ _0715_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a21o_1
XFILLER_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2335_ net139 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1217_ _0398_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1148_ P0\[20\] P0\[21\] _0903_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__mux2_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1079_ P0\[53\] P0\[54\] _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__mux2_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_23_wb_clk_i clknet_2_2__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2120_ clknet_leaf_12_wb_clk_i spm.genblk1\[24\].csa.hsum2 _0220_ VGND VGND VPWR
+ VPWR spm.genblk1\[23\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2051_ clknet_leaf_26_wb_clk_i _0338_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ net43 Y\[17\] _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__mux2_1
XFILLER_63_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1904_ clknet_leaf_23_wb_clk_i spm.genblk1\[15\].csa.hsum2 _0037_ VGND VGND VPWR
+ VPWR spm.genblk1\[14\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_187_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1835_ net131 _0602_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__and2_1
XFILLER_50_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1766_ spm.x\[19\] P0\[19\] _0669_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux2_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1697_ spm.x\[7\] P0\[7\] _0622_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__mux2_1
XFILLER_89_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ net139 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput77 net77 VGND VGND VPWR VPWR io_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_27_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput88 net88 VGND VGND VPWR VPWR io_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput99 net99 VGND VGND VPWR VPWR io_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1620_ _0596_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
XFILLER_201_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1551_ _0582_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__buf_4
XFILLER_153_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1482_ _0580_ _0581_ VGND VGND VPWR VPWR spm.genblk1\[18\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2103_ clknet_leaf_9_wb_clk_i _0390_ _0203_ VGND VGND VPWR VPWR Y\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2034_ clknet_leaf_4_wb_clk_i _0321_ _0167_ VGND VGND VPWR VPWR P0\[55\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1818_ net127 _0704_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__and2_1
XFILLER_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1749_ spm.x\[16\] P0\[16\] _0669_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__mux2_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0982_ net50 Y\[23\] _0799_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__mux2_1
XFILLER_9_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1603_ _0594_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1534_ _0587_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__inv_2
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1465_ _0541_ spm.x\[21\] _0568_ _0567_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a31o_1
XFILLER_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_230 VGND VGND VPWR VPWR SPM_example_230/HI la_data_out[44] sky130_fd_sc_hd__conb_1
XFILLER_68_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1396_ _0452_ spm.x\[31\] spm.tcmp.z VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__nand3_1
XSPM_example_241 VGND VGND VPWR VPWR SPM_example_241/HI la_data_out[55] sky130_fd_sc_hd__conb_1
XSPM_example_252 VGND VGND VPWR VPWR SPM_example_252/HI la_data_out[66] sky130_fd_sc_hd__conb_1
XFILLER_110_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_263 VGND VGND VPWR VPWR SPM_example_263/HI la_data_out[77] sky130_fd_sc_hd__conb_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSPM_example_274 VGND VGND VPWR VPWR SPM_example_274/HI la_data_out[88] sky130_fd_sc_hd__conb_1
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_285 VGND VGND VPWR VPWR SPM_example_285/HI la_data_out[99] sky130_fd_sc_hd__conb_1
XSPM_example_296 VGND VGND VPWR VPWR SPM_example_296/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2017_ clknet_leaf_25_wb_clk_i _0304_ _0150_ VGND VGND VPWR VPWR P0\[38\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ _0427_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1181_ P0\[4\] P0\[5\] _0914_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__mux2_1
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0965_ net55 Y\[28\] _0786_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__mux2_1
XFILLER_186_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1517_ _0585_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__inv_2
XFILLER_47_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1448_ spm.genblk1\[23\].csa.sc spm.genblk1\[23\].csa.y VGND VGND VPWR VPWR _0558_
+ sky130_fd_sc_hd__nor2_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1379_ _0479_ spm.x\[3\] VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__nand2_1
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1302_ spm.genblk1\[15\].csa.sc spm.genblk1\[15\].csa.y VGND VGND VPWR VPWR _0460_
+ sky130_fd_sc_hd__nor2_1
XFILLER_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1233_ _0418_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1164_ _0915_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1095_ P0\[45\] P0\[46\] _0870_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__mux2_1
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1997_ clknet_leaf_3_wb_clk_i _0284_ _0130_ VGND VGND VPWR VPWR P0\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0948_ net9 net12 net15 net16 VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__or4_1
XFILLER_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1920_ clknet_leaf_18_wb_clk_i spm.genblk1\[7\].csa.hsum2 _0053_ VGND VGND VPWR VPWR
+ spm.genblk1\[6\].csa.y sky130_fd_sc_hd__dfrtp_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1851_ _0759_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__inv_2
XFILLER_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1782_ net120 _0704_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__and2_1
XFILLER_129_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2334_ net142 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1216_ _0409_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1147_ _0906_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1078_ _0793_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__buf_4
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_8 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2050_ clknet_leaf_21_wb_clk_i _0337_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_4
XFILLER_130_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1001_ _0798_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__clkbuf_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1903_ clknet_leaf_2_wb_clk_i _0007_ _0036_ VGND VGND VPWR VPWR spm.genblk1\[16\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1834_ P0\[63\] _0611_ _0614_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__o21a_1
XFILLER_198_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1765_ _0778_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1696_ _0641_ _0642_ _0643_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a21o_1
XFILLER_171_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ net142 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_97_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_942 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput78 net78 VGND VGND VPWR VPWR io_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_153_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput89 net89 VGND VGND VPWR VPWR io_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_27_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1550_ _0588_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
XFILLER_114_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1481_ _0452_ spm.x\[18\] VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nand2_1
XFILLER_193_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2102_ clknet_leaf_7_wb_clk_i _0389_ _0202_ VGND VGND VPWR VPWR Y\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2033_ clknet_leaf_4_wb_clk_i _0320_ _0166_ VGND VGND VPWR VPWR P0\[54\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1817_ P0\[60\] _0708_ _0709_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__o21a_1
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1748_ _0684_ _0685_ _0686_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a21o_1
XFILLER_117_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1679_ net132 _0603_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__and2_1
XFILLER_85_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0981_ _0807_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1602_ _0594_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1533_ _0587_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1464_ _0568_ _0569_ VGND VGND VPWR VPWR spm.genblk1\[21\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_101_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_220 VGND VGND VPWR VPWR SPM_example_220/HI la_data_out[34] sky130_fd_sc_hd__conb_1
XFILLER_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1395_ spm.y spm.x\[31\] spm.tcmp.z VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a21o_1
XFILLER_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_231 VGND VGND VPWR VPWR SPM_example_231/HI la_data_out[45] sky130_fd_sc_hd__conb_1
XFILLER_95_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_242 VGND VGND VPWR VPWR SPM_example_242/HI la_data_out[56] sky130_fd_sc_hd__conb_1
XSPM_example_253 VGND VGND VPWR VPWR SPM_example_253/HI la_data_out[67] sky130_fd_sc_hd__conb_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_264 VGND VGND VPWR VPWR SPM_example_264/HI la_data_out[78] sky130_fd_sc_hd__conb_1
XFILLER_83_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSPM_example_275 VGND VGND VPWR VPWR SPM_example_275/HI la_data_out[89] sky130_fd_sc_hd__conb_1
XSPM_example_286 VGND VGND VPWR VPWR SPM_example_286/HI la_data_out[100] sky130_fd_sc_hd__conb_1
XSPM_example_297 VGND VGND VPWR VPWR SPM_example_297/HI la_data_out[111] sky130_fd_sc_hd__conb_1
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2016_ clknet_leaf_26_wb_clk_i _0303_ _0149_ VGND VGND VPWR VPWR P0\[37\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1180_ _0923_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0964_ _0795_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1516_ _0585_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__inv_2
XFILLER_173_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1447_ _0541_ spm.x\[24\] _0556_ _0555_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a31o_1
XFILLER_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1378_ _0510_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__nor2_1
XFILLER_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_wb_clk_i clknet_2_2__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1301_ _0455_ spm.x\[16\] _0458_ _0457_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a31o_1
XFILLER_2_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1232_ net40 spm.x\[14\] _0410_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ P0\[13\] P0\[14\] _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__mux2_1
XFILLER_93_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1094_ _0878_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ clknet_leaf_3_wb_clk_i _0283_ _0129_ VGND VGND VPWR VPWR P0\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_197_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0947_ net18 net21 net25 net23 VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__or4b_1
XFILLER_147_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1850_ _0759_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__inv_2
XFILLER_204_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1781_ P0\[53\] _0708_ _0709_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__o21a_1
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2333_ net1 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1215_ net49 spm.x\[22\] _0399_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux2_1
XFILLER_211_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1146_ P0\[21\] P0\[22\] _0903_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__mux2_1
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1077_ _0869_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1979_ clknet_leaf_17_wb_clk_i _0266_ _0112_ VGND VGND VPWR VPWR P0\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_9 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1000_ _0820_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1902_ clknet_leaf_23_wb_clk_i spm.genblk1\[16\].csa.hsum2 _0035_ VGND VGND VPWR
+ VPWR spm.genblk1\[15\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_176_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1833_ _0787_ _0754_ _0755_ _0606_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__a211o_1
XFILLER_129_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1764_ _0697_ _0698_ _0699_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a21o_1
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1695_ net135 _0603_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__and2_1
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2316_ net140 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1129_ P0\[29\] P0\[30\] _0892_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__mux2_1
XFILLER_26_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput79 net79 VGND VGND VPWR VPWR io_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_103_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1480_ _0578_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__nor2_1
XFILLER_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2101_ clknet_leaf_6_wb_clk_i _0388_ _0201_ VGND VGND VPWR VPWR Y\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2032_ clknet_leaf_4_wb_clk_i _0319_ _0165_ VGND VGND VPWR VPWR P0\[53\] sky130_fd_sc_hd__dfrtp_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1816_ Y\[28\] _0700_ _0786_ _0741_ _0605_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__a221o_1
XFILLER_163_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1747_ net113 _0657_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__and2_1
XFILLER_172_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1678_ P0\[35\] _0612_ _0615_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__o21a_1
XFILLER_172_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0980_ _0806_ Y\[25\] _0794_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__mux2_1
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1601_ _0594_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__inv_2
XFILLER_161_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1532_ _0587_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
XFILLER_114_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1463_ _0452_ spm.x\[21\] VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nand2_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_210 VGND VGND VPWR VPWR SPM_example_210/HI la_data_out[24] sky130_fd_sc_hd__conb_1
X_1394_ _0497_ spm.x\[1\] _0520_ _0519_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a31o_1
XSPM_example_221 VGND VGND VPWR VPWR SPM_example_221/HI la_data_out[35] sky130_fd_sc_hd__conb_1
XFILLER_68_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSPM_example_232 VGND VGND VPWR VPWR SPM_example_232/HI la_data_out[46] sky130_fd_sc_hd__conb_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_243 VGND VGND VPWR VPWR SPM_example_243/HI la_data_out[57] sky130_fd_sc_hd__conb_1
XFILLER_95_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_254 VGND VGND VPWR VPWR SPM_example_254/HI la_data_out[68] sky130_fd_sc_hd__conb_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_265 VGND VGND VPWR VPWR SPM_example_265/HI la_data_out[79] sky130_fd_sc_hd__conb_1
XSPM_example_276 VGND VGND VPWR VPWR SPM_example_276/HI la_data_out[90] sky130_fd_sc_hd__conb_1
XFILLER_55_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_287 VGND VGND VPWR VPWR SPM_example_287/HI la_data_out[101] sky130_fd_sc_hd__conb_1
XSPM_example_298 VGND VGND VPWR VPWR SPM_example_298/HI la_data_out[112] sky130_fd_sc_hd__conb_1
XFILLER_209_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2015_ clknet_leaf_25_wb_clk_i _0302_ _0148_ VGND VGND VPWR VPWR P0\[36\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0963_ _0792_ Y\[30\] _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__mux2_1
XFILLER_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1515_ _0585_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__inv_2
XFILLER_82_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1446_ _0556_ _0557_ VGND VGND VPWR VPWR spm.genblk1\[24\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1377_ spm.genblk1\[3\].csa.sc spm.genblk1\[3\].csa.y VGND VGND VPWR VPWR _0511_
+ sky130_fd_sc_hd__and2_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ _0458_ _0459_ VGND VGND VPWR VPWR spm.genblk1\[16\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1231_ _0417_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1162_ STATE VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ P0\[46\] P0\[47\] _0870_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__mux2_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1995_ clknet_leaf_0_wb_clk_i _0282_ _0128_ VGND VGND VPWR VPWR P0\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0946_ net10 net11 net14 net17 VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__or4_1
XFILLER_146_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1429_ _0541_ spm.x\[27\] _0544_ _0543_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a31o_1
XFILLER_56_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1780_ Y\[21\] _0700_ _0682_ _0712_ _0692_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__a221o_1
XFILLER_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2332_ net143 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1214_ _0408_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1145_ _0905_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1076_ P0\[54\] P0\[55\] _0859_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__mux2_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1978_ clknet_leaf_15_wb_clk_i nstate\[0\] _0111_ VGND VGND VPWR VPWR STATE sky130_fd_sc_hd__dfrtp_4
XFILLER_147_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ clknet_leaf_10_wb_clk_i _0008_ _0034_ VGND VGND VPWR VPWR spm.genblk1\[17\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_203_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1832_ Y\[31\] _0778_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__and2_1
XFILLER_204_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1763_ net116 _0657_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__and2_1
XFILLER_184_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1694_ P0\[38\] _0612_ _0615_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__o21a_1
XFILLER_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ net143 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1128_ _0896_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1059_ _0860_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput69 net69 VGND VGND VPWR VPWR io_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_27_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2100_ clknet_leaf_6_wb_clk_i _0387_ _0200_ VGND VGND VPWR VPWR Y\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2031_ clknet_leaf_0_wb_clk_i _0318_ _0164_ VGND VGND VPWR VPWR P0\[52\] sky130_fd_sc_hd__dfrtp_1
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1815_ spm.x\[28\] P0\[28\] _0397_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__mux2_1
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1746_ P0\[47\] _0661_ _0662_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__o21a_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1677_ Y\[3\] _0779_ _0787_ _0627_ _0606_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a221o_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1600_ _0594_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1531_ _0587_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_153_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1462_ _0566_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nor2_1
XFILLER_45_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_200 VGND VGND VPWR VPWR SPM_example_200/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_136_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1393_ _0520_ _0522_ VGND VGND VPWR VPWR spm.genblk1\[1\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_211 VGND VGND VPWR VPWR SPM_example_211/HI la_data_out[25] sky130_fd_sc_hd__conb_1
XSPM_example_222 VGND VGND VPWR VPWR SPM_example_222/HI la_data_out[36] sky130_fd_sc_hd__conb_1
XFILLER_45_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_233 VGND VGND VPWR VPWR SPM_example_233/HI la_data_out[47] sky130_fd_sc_hd__conb_1
XSPM_example_244 VGND VGND VPWR VPWR SPM_example_244/HI la_data_out[58] sky130_fd_sc_hd__conb_1
XFILLER_132_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_255 VGND VGND VPWR VPWR SPM_example_255/HI la_data_out[69] sky130_fd_sc_hd__conb_1
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_266 VGND VGND VPWR VPWR SPM_example_266/HI la_data_out[80] sky130_fd_sc_hd__conb_1
XFILLER_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_277 VGND VGND VPWR VPWR SPM_example_277/HI la_data_out[91] sky130_fd_sc_hd__conb_1
XSPM_example_288 VGND VGND VPWR VPWR SPM_example_288/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XFILLER_55_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSPM_example_299 VGND VGND VPWR VPWR SPM_example_299/HI la_data_out[113] sky130_fd_sc_hd__conb_1
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2014_ clknet_leaf_25_wb_clk_i _0301_ _0147_ VGND VGND VPWR VPWR P0\[35\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1729_ Y\[12\] _0653_ _0635_ _0670_ _0645_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__a221o_1
XFILLER_132_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0962_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__buf_4
XFILLER_159_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1514_ _0585_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__inv_2
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1445_ _0521_ spm.x\[24\] VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__nand2_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376_ spm.genblk1\[3\].csa.sc spm.genblk1\[3\].csa.y VGND VGND VPWR VPWR _0510_
+ sky130_fd_sc_hd__nor2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1230_ net41 spm.x\[15\] _0410_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_922 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_wb_clk_i clknet_2_0__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_1161_ _0913_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1092_ _0877_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1994_ clknet_leaf_0_wb_clk_i _0281_ _0127_ VGND VGND VPWR VPWR P0\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0945_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__clkbuf_4
XFILLER_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1428_ _0544_ _0545_ VGND VGND VPWR VPWR spm.genblk1\[27\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1359_ spm.genblk1\[6\].csa.sc spm.genblk1\[6\].csa.y VGND VGND VPWR VPWR _0499_
+ sky130_fd_sc_hd__and2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2331_ net141 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_152_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1213_ net50 spm.x\[23\] _0399_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1144_ P0\[22\] P0\[23\] _0903_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__mux2_1
XFILLER_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1075_ _0868_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1977_ clknet_leaf_15_wb_clk_i ncnt\[7\] _0110_ VGND VGND VPWR VPWR CNT\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ clknet_leaf_2_wb_clk_i spm.genblk1\[17\].csa.hsum2 _0033_ VGND VGND VPWR VPWR
+ spm.genblk1\[16\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1831_ spm.x\[31\] P0\[31\] _0398_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__mux2_1
XFILLER_124_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1762_ P0\[50\] _0661_ _0662_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__o21a_1
XFILLER_129_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1693_ Y\[6\] _0779_ _0635_ _0640_ _0606_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__a221o_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2314_ net142 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1127_ P0\[30\] P0\[31\] _0892_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1058_ P0\[63\] spm.csa0.sum _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ clknet_leaf_0_wb_clk_i _0317_ _0163_ VGND VGND VPWR VPWR P0\[51\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1814_ _0738_ _0739_ _0740_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a21o_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1745_ Y\[15\] _0653_ _0682_ _0683_ _0645_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a221o_1
XFILLER_89_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1676_ spm.x\[3\] P0\[3\] _0622_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux2_1
XFILLER_171_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1530_ _0587_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__inv_2
XFILLER_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1461_ spm.genblk1\[21\].csa.sc spm.genblk1\[21\].csa.y VGND VGND VPWR VPWR _0567_
+ sky130_fd_sc_hd__and2_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1392_ _0521_ spm.x\[1\] VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__nand2_1
XSPM_example_201 VGND VGND VPWR VPWR SPM_example_201/HI la_data_out[15] sky130_fd_sc_hd__conb_1
XSPM_example_212 VGND VGND VPWR VPWR SPM_example_212/HI la_data_out[26] sky130_fd_sc_hd__conb_1
XFILLER_136_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_223 VGND VGND VPWR VPWR SPM_example_223/HI la_data_out[37] sky130_fd_sc_hd__conb_1
XSPM_example_234 VGND VGND VPWR VPWR SPM_example_234/HI la_data_out[48] sky130_fd_sc_hd__conb_1
XFILLER_45_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_245 VGND VGND VPWR VPWR SPM_example_245/HI la_data_out[59] sky130_fd_sc_hd__conb_1
XFILLER_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSPM_example_256 VGND VGND VPWR VPWR SPM_example_256/HI la_data_out[70] sky130_fd_sc_hd__conb_1
XSPM_example_267 VGND VGND VPWR VPWR SPM_example_267/HI la_data_out[81] sky130_fd_sc_hd__conb_1
XSPM_example_278 VGND VGND VPWR VPWR SPM_example_278/HI la_data_out[92] sky130_fd_sc_hd__conb_1
XFILLER_94_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_289 VGND VGND VPWR VPWR SPM_example_289/HI la_data_out[103] sky130_fd_sc_hd__conb_1
X_2013_ clknet_leaf_25_wb_clk_i _0300_ _0146_ VGND VGND VPWR VPWR P0\[34\] sky130_fd_sc_hd__dfrtp_1
XFILLER_209_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1728_ spm.x\[12\] P0\[12\] _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux2_1
XFILLER_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1659_ _0769_ _0770_ _0771_ _0608_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__or4_1
XFILLER_132_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ STATE VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__buf_4
XFILLER_201_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1513_ _0585_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__inv_2
XFILLER_153_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1444_ _0554_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__nor2_1
X_1375_ _0497_ spm.x\[4\] _0508_ _0507_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a31o_1
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1160_ P0\[14\] P0\[15\] _0903_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__mux2_1
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ P0\[47\] P0\[48\] _0870_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__mux2_1
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1993_ clknet_leaf_0_wb_clk_i _0280_ _0126_ VGND VGND VPWR VPWR P0\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0944_ _0764_ _0768_ _0772_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nor4_2
XFILLER_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1427_ _0521_ spm.x\[27\] VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nand2_1
XFILLER_130_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1358_ spm.genblk1\[6\].csa.sc spm.genblk1\[6\].csa.y VGND VGND VPWR VPWR _0498_
+ sky130_fd_sc_hd__nor2_1
XFILLER_56_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1289_ _0449_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nor2_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2330_ net139 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1212_ _0407_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1143_ _0904_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1074_ P0\[55\] P0\[56\] _0859_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__mux2_1
XFILLER_81_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ clknet_leaf_15_wb_clk_i ncnt\[6\] _0109_ VGND VGND VPWR VPWR CNT\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_193_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ _0751_ _0752_ _0753_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a21o_1
XFILLER_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1761_ Y\[18\] _0653_ _0682_ _0696_ _0692_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__a221o_1
XFILLER_204_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1692_ spm.x\[6\] P0\[6\] _0622_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux2_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1007 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ net139 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1126_ _0895_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1057_ _0793_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__clkbuf_4
XFILLER_202_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1959_ clknet_leaf_3_wb_clk_i _0255_ _0092_ VGND VGND VPWR VPWR spm.x\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1813_ net126 _0704_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__and2_1
XFILLER_129_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1744_ spm.x\[15\] P0\[15\] _0669_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__mux2_1
XFILLER_129_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1675_ _0624_ _0625_ _0626_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a21o_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1109_ _0886_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__clkbuf_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2089_ clknet_leaf_0_wb_clk_i _0376_ _0189_ VGND VGND VPWR VPWR Y\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1460_ spm.genblk1\[21\].csa.sc spm.genblk1\[21\].csa.y VGND VGND VPWR VPWR _0566_
+ sky130_fd_sc_hd__nor2_1
XFILLER_45_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1391_ _0452_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__clkbuf_4
XSPM_example_202 VGND VGND VPWR VPWR SPM_example_202/HI la_data_out[16] sky130_fd_sc_hd__conb_1
XFILLER_45_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_213 VGND VGND VPWR VPWR SPM_example_213/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XSPM_example_224 VGND VGND VPWR VPWR SPM_example_224/HI la_data_out[38] sky130_fd_sc_hd__conb_1
XSPM_example_235 VGND VGND VPWR VPWR SPM_example_235/HI la_data_out[49] sky130_fd_sc_hd__conb_1
XSPM_example_246 VGND VGND VPWR VPWR SPM_example_246/HI la_data_out[60] sky130_fd_sc_hd__conb_1
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_257 VGND VGND VPWR VPWR SPM_example_257/HI la_data_out[71] sky130_fd_sc_hd__conb_1
XSPM_example_268 VGND VGND VPWR VPWR SPM_example_268/HI la_data_out[82] sky130_fd_sc_hd__conb_1
XSPM_example_279 VGND VGND VPWR VPWR SPM_example_279/HI la_data_out[93] sky130_fd_sc_hd__conb_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2012_ clknet_leaf_25_wb_clk_i _0299_ _0145_ VGND VGND VPWR VPWR P0\[33\] sky130_fd_sc_hd__dfrtp_1
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1727_ _0397_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1658_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__buf_2
XFILLER_171_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1589_ _0593_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0960_ net56 Y\[29\] _0786_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__mux2_1
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1512_ _0585_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__inv_2
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1443_ spm.genblk1\[24\].csa.sc spm.genblk1\[24\].csa.y VGND VGND VPWR VPWR _0555_
+ sky130_fd_sc_hd__and2_1
XFILLER_68_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1374_ _0508_ _0509_ VGND VGND VPWR VPWR spm.genblk1\[4\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1090_ _0876_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1992_ clknet_leaf_0_wb_clk_i _0279_ _0125_ VGND VGND VPWR VPWR P0\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0943_ _0773_ _0774_ _0775_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__or4_1
XFILLER_202_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1426_ _0542_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nor2_1
XFILLER_60_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1357_ _0497_ spm.x\[7\] _0495_ _0494_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__a31o_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1288_ spm.genblk1\[17\].csa.sc spm.genblk1\[17\].csa.y VGND VGND VPWR VPWR _0450_
+ sky130_fd_sc_hd__and2_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1211_ net51 spm.x\[24\] _0399_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux2_1
XFILLER_46_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1142_ P0\[23\] P0\[24\] _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__mux2_1
XFILLER_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1073_ _0867_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1975_ clknet_leaf_13_wb_clk_i ncnt\[5\] _0108_ VGND VGND VPWR VPWR CNT\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_105_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1409_ _0531_ _0532_ VGND VGND VPWR VPWR spm.genblk1\[30\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1760_ spm.x\[18\] P0\[18\] _0669_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux2_1
XFILLER_128_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1691_ _0637_ _0638_ _0639_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a21o_1
XFILLER_128_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2312_ net140 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1125_ P0\[31\] P0\[32\] _0892_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__mux2_1
XFILLER_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1056_ _0858_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1958_ clknet_leaf_3_wb_clk_i _0254_ _0091_ VGND VGND VPWR VPWR spm.x\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1889_ _0763_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__inv_2
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1812_ P0\[59\] _0708_ _0709_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__o21a_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1743_ _0786_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__buf_2
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1674_ net129 _0603_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__and2_1
XFILLER_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1108_ P0\[39\] P0\[40\] _0881_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__mux2_1
XFILLER_96_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2088_ clknet_leaf_28_wb_clk_i _0375_ _0188_ VGND VGND VPWR VPWR Y\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1039_ net62 Y\[5\] _0798_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__mux2_1
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ _0518_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__nor2_1
XFILLER_171_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_203 VGND VGND VPWR VPWR SPM_example_203/HI la_data_out[17] sky130_fd_sc_hd__conb_1
XSPM_example_214 VGND VGND VPWR VPWR SPM_example_214/HI la_data_out[28] sky130_fd_sc_hd__conb_1
XFILLER_45_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_225 VGND VGND VPWR VPWR SPM_example_225/HI la_data_out[39] sky130_fd_sc_hd__conb_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_236 VGND VGND VPWR VPWR SPM_example_236/HI la_data_out[50] sky130_fd_sc_hd__conb_1
XSPM_example_247 VGND VGND VPWR VPWR SPM_example_247/HI la_data_out[61] sky130_fd_sc_hd__conb_1
XSPM_example_258 VGND VGND VPWR VPWR SPM_example_258/HI la_data_out[72] sky130_fd_sc_hd__conb_1
XFILLER_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_269 VGND VGND VPWR VPWR SPM_example_269/HI la_data_out[83] sky130_fd_sc_hd__conb_1
XFILLER_208_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ clknet_leaf_25_wb_clk_i _0298_ _0144_ VGND VGND VPWR VPWR P0\[32\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1726_ _0666_ _0667_ _0668_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a21o_1
XFILLER_208_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1657_ _0764_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or2_2
XFILLER_208_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1588_ _0593_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1511_ _0585_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__inv_2
XFILLER_182_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1442_ spm.genblk1\[24\].csa.sc spm.genblk1\[24\].csa.y VGND VGND VPWR VPWR _0554_
+ sky130_fd_sc_hd__nor2_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1373_ _0479_ spm.x\[4\] VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__nand2_1
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1082 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1709_ spm.x\[9\] P0\[9\] _0622_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux2_1
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1991_ clknet_leaf_28_wb_clk_i _0278_ _0124_ VGND VGND VPWR VPWR P0\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0942_ net26 net25 net23 net22 VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__or4bb_1
XFILLER_140_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1425_ spm.genblk1\[27\].csa.sc spm.genblk1\[27\].csa.y VGND VGND VPWR VPWR _0543_
+ sky130_fd_sc_hd__and2_1
XFILLER_130_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1356_ _0453_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1287_ spm.genblk1\[17\].csa.sc spm.genblk1\[17\].csa.y VGND VGND VPWR VPWR _0449_
+ sky130_fd_sc_hd__nor2_1
XFILLER_3_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1210_ _0406_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1141_ STATE VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_120_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1072_ P0\[56\] P0\[57\] _0859_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__mux2_1
XFILLER_207_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ clknet_leaf_13_wb_clk_i ncnt\[4\] _0107_ VGND VGND VPWR VPWR CNT\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1408_ _0521_ spm.x\[30\] VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__nand2_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1339_ spm.genblk1\[9\].csa.sc spm.genblk1\[10\].csa.sum VGND VGND VPWR VPWR _0485_
+ sky130_fd_sc_hd__nor2_1
XFILLER_186_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1690_ net134 _0603_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__and2_1
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2311_ net143 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_152_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1124_ _0894_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1055_ _0857_ Y\[1\] _0839_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__mux2_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1957_ clknet_leaf_3_wb_clk_i _0253_ _0090_ VGND VGND VPWR VPWR spm.x\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1888_ net142 VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__buf_4
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _0787_ _0736_ _0737_ _0606_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a211o_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1742_ _0679_ _0680_ _0681_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a21o_1
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1673_ P0\[34\] _0612_ _0615_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__o21a_1
XFILLER_144_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1107_ _0885_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2087_ clknet_leaf_24_wb_clk_i _0374_ _0187_ VGND VGND VPWR VPWR Y\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1038_ _0846_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_204 VGND VGND VPWR VPWR SPM_example_204/HI la_data_out[18] sky130_fd_sc_hd__conb_1
XFILLER_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_215 VGND VGND VPWR VPWR SPM_example_215/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_110_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_226 VGND VGND VPWR VPWR SPM_example_226/HI la_data_out[40] sky130_fd_sc_hd__conb_1
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_237 VGND VGND VPWR VPWR SPM_example_237/HI la_data_out[51] sky130_fd_sc_hd__conb_1
XSPM_example_248 VGND VGND VPWR VPWR SPM_example_248/HI la_data_out[62] sky130_fd_sc_hd__conb_1
XFILLER_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_259 VGND VGND VPWR VPWR SPM_example_259/HI la_data_out[73] sky130_fd_sc_hd__conb_1
X_2010_ clknet_leaf_24_wb_clk_i _0297_ _0143_ VGND VGND VPWR VPWR P0\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1725_ net109 _0657_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and2_1
XFILLER_145_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1656_ _0929_ _0608_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or3_1
XFILLER_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1587_ _0593_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1510_ _0585_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__inv_2
XFILLER_99_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1441_ _0541_ spm.x\[25\] _0552_ _0551_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a31o_1
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1372_ _0506_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__nor2_1
XFILLER_68_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1094 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1708_ _0778_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__clkbuf_4
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1639_ _0597_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__inv_2
XFILLER_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1990_ clknet_leaf_1_wb_clk_i _0277_ _0123_ VGND VGND VPWR VPWR P0\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ net19 net18 net21 net20 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__or4_1
XFILLER_201_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1424_ spm.genblk1\[27\].csa.sc spm.genblk1\[27\].csa.y VGND VGND VPWR VPWR _0542_
+ sky130_fd_sc_hd__nor2_1
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1355_ _0495_ _0496_ VGND VGND VPWR VPWR spm.genblk1\[7\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_60_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1286_ CNT\[7\] _0446_ _0448_ VGND VGND VPWR VPWR ncnt\[7\] sky130_fd_sc_hd__a21oi_1
XFILLER_49_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1140_ _0902_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1071_ _0866_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ clknet_leaf_14_wb_clk_i ncnt\[3\] _0106_ VGND VGND VPWR VPWR CNT\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_105_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1407_ _0529_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1338_ _0455_ spm.x\[10\] _0483_ _0482_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a31o_1
XFILLER_112_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1269_ CNT\[1\] CNT\[0\] _0437_ VGND VGND VPWR VPWR ncnt\[1\] sky130_fd_sc_hd__a21oi_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2310_ net143 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1123_ P0\[32\] P0\[33\] _0892_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__mux2_1
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1054_ net35 spm.y _0798_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__mux2_1
XFILLER_202_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1956_ clknet_leaf_2_wb_clk_i _0252_ _0089_ VGND VGND VPWR VPWR spm.x\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1887_ _0762_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__inv_2
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1810_ Y\[27\] _0778_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and2_1
XFILLER_54_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1741_ net112 _0657_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and2_1
XFILLER_89_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1672_ Y\[2\] _0779_ _0787_ _0623_ _0606_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a221o_1
XFILLER_183_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1106_ P0\[40\] P0\[41\] _0881_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__mux2_1
XFILLER_199_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2086_ clknet_leaf_23_wb_clk_i _0373_ _0186_ VGND VGND VPWR VPWR Y\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1037_ _0845_ Y\[7\] _0839_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__mux2_1
XFILLER_22_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1939_ clknet_leaf_16_wb_clk_i _0235_ _0072_ VGND VGND VPWR VPWR spm.x\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_205 VGND VGND VPWR VPWR SPM_example_205/HI la_data_out[19] sky130_fd_sc_hd__conb_1
XSPM_example_216 VGND VGND VPWR VPWR SPM_example_216/HI la_data_out[30] sky130_fd_sc_hd__conb_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_227 VGND VGND VPWR VPWR SPM_example_227/HI la_data_out[41] sky130_fd_sc_hd__conb_1
XFILLER_110_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_238 VGND VGND VPWR VPWR SPM_example_238/HI la_data_out[52] sky130_fd_sc_hd__conb_1
XSPM_example_249 VGND VGND VPWR VPWR SPM_example_249/HI la_data_out[63] sky130_fd_sc_hd__conb_1
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1724_ P0\[43\] _0661_ _0662_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__o21a_1
XFILLER_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1655_ net68 _0599_ _0770_ _0771_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__or4_1
XFILLER_208_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1586_ _0593_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
XFILLER_99_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2069_ clknet_leaf_5_wb_clk_i _0356_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_4
XFILLER_156_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1440_ _0552_ _0553_ VGND VGND VPWR VPWR spm.genblk1\[25\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_175_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1371_ spm.genblk1\[4\].csa.sc spm.genblk1\[4\].csa.y VGND VGND VPWR VPWR _0507_
+ sky130_fd_sc_hd__and2_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1707_ _0650_ _0651_ _0652_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a21o_1
XFILLER_160_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1638_ _0597_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__inv_2
XFILLER_8_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1569_ _0590_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
XFILLER_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ net10 net9 net12 net11 VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__or4_1
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1423_ _0541_ spm.x\[28\] _0539_ _0538_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a31o_1
XFILLER_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1354_ _0479_ spm.x\[7\] VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__nand2_1
XFILLER_205_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1285_ CNT\[7\] _0446_ _0788_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__o21ai_1
XFILLER_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clknet_2_3__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1070_ P0\[57\] P0\[58\] _0859_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__mux2_1
XFILLER_207_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1972_ clknet_leaf_14_wb_clk_i ncnt\[2\] _0105_ VGND VGND VPWR VPWR CNT\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1406_ spm.genblk1\[30\].csa.sc spm.genblk1\[30\].csa.y VGND VGND VPWR VPWR _0530_
+ sky130_fd_sc_hd__and2_1
XFILLER_151_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1337_ _0483_ _0484_ VGND VGND VPWR VPWR spm.genblk1\[10\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_25_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1268_ CNT\[1\] CNT\[0\] _0788_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1199_ net58 spm.x\[30\] _0399_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux2_1
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1122_ _0893_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1053_ _0856_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1955_ clknet_leaf_2_wb_clk_i _0251_ _0088_ VGND VGND VPWR VPWR spm.x\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1886_ _0762_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__inv_2
XFILLER_190_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_60 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1740_ P0\[46\] _0661_ _0662_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__o21a_1
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1671_ spm.x\[2\] P0\[2\] _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1105_ _0884_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2085_ clknet_leaf_23_wb_clk_i _0372_ _0185_ VGND VGND VPWR VPWR Y\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1036_ net63 Y\[6\] _0798_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__mux2_1
XFILLER_62_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1938_ clknet_leaf_15_wb_clk_i _0234_ _0071_ VGND VGND VPWR VPWR spm.x\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_120_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1869_ _0761_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__inv_2
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_206 VGND VGND VPWR VPWR SPM_example_206/HI la_data_out[20] sky130_fd_sc_hd__conb_1
XSPM_example_217 VGND VGND VPWR VPWR SPM_example_217/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSPM_example_228 VGND VGND VPWR VPWR SPM_example_228/HI la_data_out[42] sky130_fd_sc_hd__conb_1
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_239 VGND VGND VPWR VPWR SPM_example_239/HI la_data_out[53] sky130_fd_sc_hd__conb_1
XFILLER_209_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1723_ Y\[11\] _0653_ _0635_ _0665_ _0645_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__a221o_1
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1654_ _0773_ _0774_ _0775_ _0776_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or4_1
XFILLER_99_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1585_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__buf_4
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2068_ clknet_leaf_4_wb_clk_i _0355_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_2
XFILLER_82_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1019_ _0833_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1370_ spm.genblk1\[4\].csa.sc spm.genblk1\[4\].csa.y VGND VGND VPWR VPWR _0506_
+ sky130_fd_sc_hd__nor2_1
XFILLER_96_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1706_ net137 _0603_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__and2_1
XFILLER_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1637_ _0597_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__inv_2
XFILLER_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1568_ _0590_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1499_ _0584_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1422_ _0453_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1353_ _0493_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nor2_1
XFILLER_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1284_ _0436_ _0446_ _0447_ VGND VGND VPWR VPWR ncnt\[6\] sky130_fd_sc_hd__nor3_1
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0999_ _0819_ Y\[19\] _0817_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__mux2_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1971_ clknet_leaf_14_wb_clk_i ncnt\[1\] _0104_ VGND VGND VPWR VPWR CNT\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1405_ spm.genblk1\[30\].csa.sc spm.genblk1\[30\].csa.y VGND VGND VPWR VPWR _0529_
+ sky130_fd_sc_hd__nor2_1
XFILLER_190_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1336_ _0479_ spm.x\[10\] VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nand2_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 wb_rst_i VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_6
XFILLER_151_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1267_ CNT\[0\] _0436_ VGND VGND VPWR VPWR ncnt\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_37_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1198_ _0400_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1121_ P0\[33\] P0\[34\] _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__mux2_1
XFILLER_19_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1052_ _0855_ Y\[2\] _0839_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__mux2_1
XFILLER_207_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1954_ clknet_leaf_1_wb_clk_i _0250_ _0087_ VGND VGND VPWR VPWR spm.x\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1885_ _0762_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__inv_2
XFILLER_175_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1319_ _0455_ spm.x\[13\] _0470_ _0469_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a31o_1
XFILLER_186_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_50 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_61 net142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1670_ _0397_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__clkbuf_4
XFILLER_176_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1104_ P0\[41\] P0\[42\] _0881_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__mux2_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2084_ clknet_leaf_23_wb_clk_i _0371_ _0184_ VGND VGND VPWR VPWR Y\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1035_ _0844_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1937_ clknet_leaf_15_wb_clk_i _0000_ _0070_ VGND VGND VPWR VPWR spm.csa0.sc sky130_fd_sc_hd__dfrtp_1
XFILLER_175_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1868_ _0761_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__inv_2
XFILLER_200_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1799_ spm.x\[25\] P0\[25\] _0397_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__mux2_1
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_199_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_207 VGND VGND VPWR VPWR SPM_example_207/HI la_data_out[21] sky130_fd_sc_hd__conb_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_218 VGND VGND VPWR VPWR SPM_example_218/HI la_data_out[32] sky130_fd_sc_hd__conb_1
XSPM_example_229 VGND VGND VPWR VPWR SPM_example_229/HI la_data_out[43] sky130_fd_sc_hd__conb_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1722_ spm.x\[11\] P0\[11\] _0622_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__mux2_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1653_ _0452_ _0779_ _0787_ _0604_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__a221o_1
XFILLER_176_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1584_ net142 VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__buf_4
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2067_ clknet_leaf_4_wb_clk_i _0354_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_2
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1018_ _0832_ Y\[13\] _0817_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__mux2_1
XFILLER_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1705_ P0\[40\] _0612_ _0615_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o21a_1
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1636_ _0597_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__inv_2
XFILLER_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1567_ _0590_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
XFILLER_113_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1498_ _0584_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XFILLER_87_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2119_ clknet_leaf_7_wb_clk_i _0017_ _0219_ VGND VGND VPWR VPWR spm.genblk1\[25\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1421_ _0539_ _0540_ VGND VGND VPWR VPWR spm.genblk1\[28\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1352_ spm.genblk1\[7\].csa.sc spm.genblk1\[7\].csa.y VGND VGND VPWR VPWR _0494_
+ sky130_fd_sc_hd__and2_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1283_ CNT\[5\] _0443_ CNT\[6\] VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a21oi_1
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0998_ net44 Y\[18\] _0799_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_wb_clk_i clknet_2_2__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1619_ _0596_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__inv_2
XFILLER_121_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ clknet_leaf_15_wb_clk_i ncnt\[0\] _0103_ VGND VGND VPWR VPWR CNT\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1404_ _0497_ spm.x\[0\] _0527_ _0526_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a31o_1
XFILLER_151_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1335_ _0481_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nor2_1
XFILLER_151_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 wbs_adr_i[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1266_ _0788_ _0787_ _0436_ VGND VGND VPWR VPWR nstate\[0\] sky130_fd_sc_hd__o21ai_1
XFILLER_37_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1197_ net59 spm.x\[31\] _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
XFILLER_188_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1120_ STATE VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__buf_4
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1051_ net46 Y\[1\] _0798_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1953_ clknet_leaf_1_wb_clk_i _0249_ _0086_ VGND VGND VPWR VPWR spm.x\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1884_ _0762_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__inv_2
XFILLER_174_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1318_ _0470_ _0471_ VGND VGND VPWR VPWR spm.genblk1\[13\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_116_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1249_ net63 spm.x\[6\] _0421_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_40 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_51 net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_62 net143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1103_ _0883_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2083_ clknet_leaf_24_wb_clk_i _0370_ _0183_ VGND VGND VPWR VPWR Y\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1034_ _0843_ Y\[8\] _0839_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__mux2_1
XFILLER_207_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1936_ clknet_leaf_15_wb_clk_i spm.csa0.hsum2 _0069_ VGND VGND VPWR VPWR spm.csa0.sum
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1867_ _0761_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__inv_2
XFILLER_135_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput60 wbs_dat_i[3] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_190_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1798_ _0725_ _0726_ _0727_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__a21o_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_208 VGND VGND VPWR VPWR SPM_example_208/HI la_data_out[22] sky130_fd_sc_hd__conb_1
XFILLER_164_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_219 VGND VGND VPWR VPWR SPM_example_219/HI la_data_out[33] sky130_fd_sc_hd__conb_1
XFILLER_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1721_ _0660_ _0663_ _0664_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__a21o_1
XFILLER_172_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1652_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1583_ _0591_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2066_ clknet_leaf_6_wb_clk_i _0353_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_4
XFILLER_208_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1017_ net38 Y\[12\] _0821_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__mux2_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1919_ clknet_leaf_17_wb_clk_i _0029_ _0052_ VGND VGND VPWR VPWR spm.genblk1\[8\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_191_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1704_ Y\[8\] _0779_ _0635_ _0649_ _0645_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__a221o_1
XFILLER_173_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635_ _0597_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
XFILLER_144_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1566_ _0590_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
XFILLER_28_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1497_ _0584_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
XFILLER_87_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2118_ clknet_leaf_7_wb_clk_i spm.genblk1\[25\].csa.hsum2 _0218_ VGND VGND VPWR VPWR
+ spm.genblk1\[24\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ clknet_leaf_26_wb_clk_i _0336_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_4
XFILLER_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1420_ _0521_ spm.x\[28\] VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand2_1
XFILLER_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1351_ spm.genblk1\[7\].csa.sc spm.genblk1\[7\].csa.y VGND VGND VPWR VPWR _0493_
+ sky130_fd_sc_hd__nor2_1
XFILLER_110_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1282_ CNT\[5\] CNT\[6\] _0443_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__and3_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0997_ _0818_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1618_ _0592_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__buf_4
XFILLER_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1549_ _0588_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
XFILLER_8_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_971 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1403_ _0527_ _0528_ VGND VGND VPWR VPWR spm.csa0.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_142_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1334_ spm.genblk1\[10\].csa.sc spm.genblk1\[10\].csa.y VGND VGND VPWR VPWR _0482_
+ sky130_fd_sc_hd__and2_1
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1265_ _0434_ _0435_ _0788_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__o21ai_1
Xinput3 wbs_adr_i[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1196_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__buf_4
XFILLER_149_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1050_ _0854_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ clknet_leaf_1_wb_clk_i _0248_ _0085_ VGND VGND VPWR VPWR spm.x\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1883_ _0762_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__inv_2
XFILLER_31_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1317_ _0453_ spm.x\[13\] VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_42_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1248_ _0426_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1179_ P0\[5\] P0\[6\] _0914_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__mux2_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_30 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1102_ P0\[42\] P0\[43\] _0881_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__mux2_1
X_2082_ clknet_leaf_25_wb_clk_i _0369_ _0182_ VGND VGND VPWR VPWR Y\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1033_ net64 Y\[7\] _0798_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__mux2_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1935_ clknet_leaf_15_wb_clk_i _0032_ _0068_ VGND VGND VPWR VPWR spm.tcmp.z sky130_fd_sc_hd__dfrtp_1
XFILLER_175_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1866_ _0592_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__buf_4
XFILLER_174_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput50 wbs_dat_i[23] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_135_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput61 wbs_dat_i[4] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1797_ net123 _0704_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__and2_1
XFILLER_190_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_209 VGND VGND VPWR VPWR SPM_example_209/HI la_data_out[23] sky130_fd_sc_hd__conb_1
XFILLER_48_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1720_ net108 _0657_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and2_1
XFILLER_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1651_ _0764_ _0601_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__nor2_2
XFILLER_176_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1582_ _0591_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2065_ clknet_leaf_4_wb_clk_i _0352_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1016_ _0831_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_wb_clk_i clknet_2_3__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1918_ clknet_leaf_18_wb_clk_i spm.genblk1\[8\].csa.hsum2 _0051_ VGND VGND VPWR VPWR
+ spm.genblk1\[7\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_120_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1849_ _0759_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__inv_2
XFILLER_194_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1703_ spm.x\[8\] P0\[8\] _0622_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1634_ _0597_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__inv_2
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1565_ _0590_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
XFILLER_98_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1496_ _0582_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__buf_4
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2117_ clknet_leaf_8_wb_clk_i _0018_ _0217_ VGND VGND VPWR VPWR spm.genblk1\[26\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2048_ clknet_leaf_26_wb_clk_i _0335_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_2
XFILLER_82_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1350_ _0455_ spm.x\[8\] _0491_ _0490_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a31o_1
XFILLER_110_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1281_ CNT\[5\] _0443_ _0445_ VGND VGND VPWR VPWR ncnt\[5\] sky130_fd_sc_hd__a21oi_1
XFILLER_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0996_ _0816_ Y\[20\] _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1617_ _0595_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__inv_2
XFILLER_99_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1548_ _0588_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
XFILLER_99_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1479_ spm.genblk1\[18\].csa.sc spm.genblk1\[18\].csa.y VGND VGND VPWR VPWR _0579_
+ sky130_fd_sc_hd__and2_1
XFILLER_80_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1402_ _0521_ spm.x\[0\] VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__nand2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1333_ spm.genblk1\[10\].csa.sc spm.genblk1\[10\].csa.y VGND VGND VPWR VPWR _0481_
+ sky130_fd_sc_hd__nor2_1
XFILLER_110_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1264_ CNT\[1\] CNT\[0\] CNT\[3\] CNT\[2\] VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or4_1
Xinput4 wbs_adr_i[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
XFILLER_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1195_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__buf_4
XFILLER_65_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0979_ net51 Y\[24\] _0799_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__mux2_1
XFILLER_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ clknet_leaf_1_wb_clk_i _0247_ _0084_ VGND VGND VPWR VPWR spm.x\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1882_ _0762_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__inv_2
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1316_ _0468_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__nor2_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1247_ net64 spm.x\[7\] _0421_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1178_ _0922_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_20 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_31 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_42 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_64 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1101_ _0882_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__clkbuf_1
X_2081_ clknet_leaf_25_wb_clk_i _0368_ _0181_ VGND VGND VPWR VPWR Y\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1032_ _0842_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1934_ clknet_leaf_15_wb_clk_i _0031_ _0067_ VGND VGND VPWR VPWR spm.genblk1\[30\].csa.y
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_174_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1865_ _0760_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__inv_2
Xinput40 wbs_dat_i[14] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_4
XFILLER_174_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 wbs_dat_i[24] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
Xinput62 wbs_dat_i[5] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
X_1796_ P0\[56\] _0708_ _0709_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__o21a_1
XFILLER_122_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1650_ spm.x\[0\] P0\[0\] _0398_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux2_1
XFILLER_172_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1581_ _0591_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_99_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2133_ clknet_leaf_16_wb_clk_i _0009_ _0233_ VGND VGND VPWR VPWR spm.genblk1\[18\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2064_ clknet_leaf_4_wb_clk_i _0351_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_2
XFILLER_187_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1015_ _0830_ Y\[14\] _0817_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__mux2_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1917_ clknet_leaf_17_wb_clk_i _0030_ _0050_ VGND VGND VPWR VPWR spm.genblk1\[9\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1848_ _0759_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__inv_2
XFILLER_190_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1779_ spm.x\[21\] P0\[21\] _0669_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__mux2_1
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1702_ _0646_ _0647_ _0648_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a21o_1
XFILLER_157_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1633_ _0597_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__inv_2
XFILLER_133_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1564_ _0590_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
XFILLER_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1495_ _0583_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
XFILLER_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2116_ clknet_leaf_7_wb_clk_i spm.genblk1\[26\].csa.hsum2 _0216_ VGND VGND VPWR VPWR
+ spm.genblk1\[25\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2047_ clknet_leaf_25_wb_clk_i _0334_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_2
XFILLER_78_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clknet_2_0__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1280_ CNT\[5\] _0443_ _0788_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0995_ _0793_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__buf_4
XFILLER_121_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1616_ _0595_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__inv_2
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1547_ _0588_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1478_ spm.genblk1\[18\].csa.sc spm.genblk1\[18\].csa.y VGND VGND VPWR VPWR _0578_
+ sky130_fd_sc_hd__nor2_1
XFILLER_41_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1401_ _0525_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__nor2_1
XFILLER_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1332_ _0455_ spm.x\[11\] _0478_ _0477_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a31o_1
XFILLER_25_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1263_ CNT\[5\] CNT\[4\] CNT\[7\] CNT\[6\] VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__or4b_1
XFILLER_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 wbs_adr_i[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1194_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__buf_4
XFILLER_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0978_ _0805_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_190 VGND VGND VPWR VPWR SPM_example_190/HI la_data_out[4] sky130_fd_sc_hd__conb_1
XFILLER_167_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ clknet_leaf_1_wb_clk_i _0246_ _0083_ VGND VGND VPWR VPWR spm.x\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1881_ _0762_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__inv_2
XFILLER_187_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1315_ spm.genblk1\[13\].csa.sc spm.genblk1\[13\].csa.y VGND VGND VPWR VPWR _0469_
+ sky130_fd_sc_hd__and2_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1246_ _0425_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1177_ P0\[6\] P0\[7\] _0914_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__mux2_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_32 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_43 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1100_ P0\[43\] P0\[44\] _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__mux2_1
X_2080_ clknet_leaf_21_wb_clk_i _0367_ _0180_ VGND VGND VPWR VPWR Y\[4\] sky130_fd_sc_hd__dfrtp_1
X_1031_ _0841_ Y\[9\] _0839_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__mux2_1
XFILLER_34_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ clknet_leaf_15_wb_clk_i _0011_ _0066_ VGND VGND VPWR VPWR spm.genblk1\[1\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1864_ _0760_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__inv_2
XFILLER_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 wbs_adr_i[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 wbs_dat_i[15] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xinput52 wbs_dat_i[25] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
XFILLER_116_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1795_ Y\[24\] _0700_ _0682_ _0724_ _0692_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a221o_1
Xinput63 wbs_dat_i[6] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
XFILLER_190_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1229_ _0416_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1580_ _0591_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2132_ clknet_leaf_16_wb_clk_i spm.genblk1\[18\].csa.hsum2 _0232_ VGND VGND VPWR
+ VPWR spm.genblk1\[17\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2063_ clknet_leaf_28_wb_clk_i _0350_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_4
XFILLER_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1014_ net39 Y\[13\] _0821_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__mux2_1
XFILLER_207_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1916_ clknet_leaf_17_wb_clk_i spm.genblk1\[9\].csa.hsum2 _0049_ VGND VGND VPWR VPWR
+ spm.genblk1\[8\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1847_ _0759_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__inv_2
XFILLER_135_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i clknet_2_0__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1778_ _0707_ _0710_ _0711_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a21o_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1701_ net136 _0603_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__and2_1
XFILLER_172_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1632_ _0597_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__inv_2
XFILLER_67_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1563_ _0590_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
XFILLER_99_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1494_ _0583_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2115_ clknet_leaf_12_wb_clk_i _0019_ _0215_ VGND VGND VPWR VPWR spm.genblk1\[27\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2046_ clknet_leaf_21_wb_clk_i _0333_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_1
XFILLER_208_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0994_ net45 Y\[19\] _0799_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__mux2_1
XFILLER_164_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1615_ _0595_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__inv_2
XFILLER_133_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1546_ _0588_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1477_ _0541_ spm.x\[19\] _0576_ _0575_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a31o_1
XFILLER_115_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2029_ clknet_leaf_28_wb_clk_i _0316_ _0162_ VGND VGND VPWR VPWR P0\[50\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ spm.csa0.sc spm.csa0.y VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__and2_1
XFILLER_155_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1331_ _0478_ _0480_ VGND VGND VPWR VPWR spm.genblk1\[11\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1262_ _0433_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput6 wbs_adr_i[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1193_ _0929_ _0772_ _0784_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__or4_1
XFILLER_188_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ _0804_ Y\[26\] _0794_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__mux2_1
XFILLER_118_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1529_ _0582_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__buf_4
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_180 VGND VGND VPWR VPWR SPM_example_180/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_191 VGND VGND VPWR VPWR SPM_example_191/HI la_data_out[5] sky130_fd_sc_hd__conb_1
XFILLER_210_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1880_ _0762_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__inv_2
XFILLER_186_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1314_ spm.genblk1\[13\].csa.sc spm.genblk1\[13\].csa.y VGND VGND VPWR VPWR _0468_
+ sky130_fd_sc_hd__nor2_1
XFILLER_97_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1245_ net65 spm.x\[8\] _0421_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1176_ _0921_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_44 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_55 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_66 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1030_ net65 Y\[8\] _0821_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__mux2_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_980 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ clknet_leaf_15_wb_clk_i spm.genblk1\[1\].csa.hsum2 _0065_ VGND VGND VPWR VPWR
+ spm.csa0.y sky130_fd_sc_hd__dfrtp_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1863_ _0760_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__inv_2
XFILLER_147_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 wbs_adr_i[26] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_4
Xinput31 wbs_adr_i[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 wbs_dat_i[16] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
X_1794_ spm.x\[24\] P0\[24\] _0397_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__mux2_1
Xinput53 wbs_dat_i[26] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
XFILLER_116_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput64 wbs_dat_i[7] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_4
XFILLER_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_1228_ net42 spm.x\[16\] _0410_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_26_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1159_ _0912_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2131_ clknet_leaf_10_wb_clk_i _0010_ _0231_ VGND VGND VPWR VPWR spm.genblk1\[19\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2062_ clknet_leaf_27_wb_clk_i _0349_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1013_ _0829_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1915_ clknet_leaf_17_wb_clk_i _0001_ _0048_ VGND VGND VPWR VPWR spm.genblk1\[10\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1846_ _0759_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__inv_2
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1777_ net119 _0704_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__and2_1
XFILLER_190_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2329_ net139 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1700_ P0\[39\] _0612_ _0615_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__o21a_1
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1631_ _0597_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
XFILLER_32_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1562_ _0582_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__buf_4
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1493_ _0583_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
XFILLER_67_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2114_ clknet_leaf_12_wb_clk_i spm.genblk1\[27\].csa.hsum2 _0214_ VGND VGND VPWR
+ VPWR spm.genblk1\[26\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_67_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2045_ clknet_leaf_21_wb_clk_i _0332_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1829_ net130 _0602_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__and2_1
XFILLER_117_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0993_ _0815_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1614_ _0595_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__inv_2
XFILLER_172_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1545_ _0588_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
XFILLER_125_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1476_ _0576_ _0577_ VGND VGND VPWR VPWR spm.genblk1\[19\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_141_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2028_ clknet_leaf_27_wb_clk_i _0315_ _0161_ VGND VGND VPWR VPWR P0\[49\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1330_ _0479_ spm.x\[11\] VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nand2_1
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1261_ net35 spm.x\[0\] _0398_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_1
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 wbs_adr_i[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1192_ net27 net24 VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__or2_1
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0976_ net52 Y\[25\] _0799_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__mux2_1
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1528_ _0586_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
XFILLER_82_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1459_ _0541_ spm.x\[22\] _0564_ _0563_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__a31o_1
XFILLER_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_170 VGND VGND VPWR VPWR SPM_example_170/HI io_out[25] sky130_fd_sc_hd__conb_1
XFILLER_132_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_181 VGND VGND VPWR VPWR SPM_example_181/HI io_out[36] sky130_fd_sc_hd__conb_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_192 VGND VGND VPWR VPWR SPM_example_192/HI la_data_out[6] sky130_fd_sc_hd__conb_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1313_ _0455_ spm.x\[14\] _0466_ _0465_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a31o_1
XFILLER_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1244_ _0424_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1175_ P0\[7\] P0\[8\] _0914_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_wb_clk_i clknet_2_2__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_23 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_34 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_67 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0959_ _0791_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_47_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1931_ clknet_leaf_17_wb_clk_i _0022_ _0064_ VGND VGND VPWR VPWR spm.genblk1\[2\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1862_ _0760_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__inv_2
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput10 wbs_adr_i[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
Xinput21 wbs_adr_i[27] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
XFILLER_163_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput32 wbs_adr_i[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
X_1793_ _0721_ _0722_ _0723_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a21o_1
Xinput43 wbs_dat_i[17] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput54 wbs_dat_i[27] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_4
Xinput65 wbs_dat_i[8] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
XFILLER_116_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1227_ _0415_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1158_ P0\[15\] P0\[16\] _0903_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__mux2_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1089_ P0\[48\] P0\[49\] _0870_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2130_ clknet_leaf_16_wb_clk_i spm.genblk1\[19\].csa.hsum2 _0230_ VGND VGND VPWR
+ VPWR spm.genblk1\[18\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2061_ clknet_leaf_27_wb_clk_i _0348_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_2
XFILLER_82_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1012_ _0828_ Y\[15\] _0817_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__mux2_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1914_ clknet_leaf_17_wb_clk_i spm.genblk1\[10\].csa.hsum2 _0047_ VGND VGND VPWR
+ VPWR spm.genblk1\[10\].csa.sum sky130_fd_sc_hd__dfrtp_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1845_ _0759_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__inv_2
XFILLER_163_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1776_ P0\[52\] _0708_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__o21a_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2328_ net143 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1630_ _0597_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__inv_2
XFILLER_67_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1561_ _0589_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1492_ _0583_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_2
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2113_ clknet_leaf_11_wb_clk_i _0020_ _0213_ VGND VGND VPWR VPWR spm.genblk1\[28\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2044_ clknet_leaf_21_wb_clk_i _0331_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_4
XFILLER_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1828_ P0\[62\] _0611_ _0614_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__o21a_1
XFILLER_190_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1759_ _0693_ _0694_ _0695_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a21o_1
XFILLER_190_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0992_ _0814_ Y\[21\] _0794_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__mux2_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1613_ _0595_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
XFILLER_172_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1544_ _0588_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
XFILLER_119_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1475_ _0452_ spm.x\[19\] VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__nand2_1
XFILLER_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2027_ clknet_leaf_27_wb_clk_i _0314_ _0160_ VGND VGND VPWR VPWR P0\[48\] sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1260_ _0432_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_2_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1191_ _0765_ _0766_ _0767_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__or3_2
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 wbs_adr_i[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0975_ _0803_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1527_ _0586_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
XFILLER_141_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1458_ _0564_ _0565_ VGND VGND VPWR VPWR spm.genblk1\[22\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_210_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_160 VGND VGND VPWR VPWR SPM_example_160/HI io_out[15] sky130_fd_sc_hd__conb_1
XFILLER_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_171 VGND VGND VPWR VPWR SPM_example_171/HI io_out[26] sky130_fd_sc_hd__conb_1
X_1389_ spm.genblk1\[1\].csa.sc spm.genblk1\[1\].csa.y VGND VGND VPWR VPWR _0519_
+ sky130_fd_sc_hd__and2_1
XFILLER_110_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_182 VGND VGND VPWR VPWR SPM_example_182/HI io_out[37] sky130_fd_sc_hd__conb_1
XFILLER_132_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_193 VGND VGND VPWR VPWR SPM_example_193/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1312_ _0466_ _0467_ VGND VGND VPWR VPWR spm.genblk1\[14\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1243_ net66 spm.x\[9\] _0421_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
XFILLER_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1174_ _0920_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_13 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_24 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_35 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_46 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_68 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0958_ _0790_ Y\[31\] _0788_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__mux2_1
XFILLER_118_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput120 net120 VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput131 net131 VGND VGND VPWR VPWR wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ clknet_leaf_17_wb_clk_i spm.genblk1\[2\].csa.hsum2 _0063_ VGND VGND VPWR VPWR
+ spm.genblk1\[1\].csa.y sky130_fd_sc_hd__dfrtp_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1861_ _0760_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__inv_2
XFILLER_147_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput11 wbs_adr_i[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput22 wbs_adr_i[28] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1792_ net122 _0704_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__and2_1
Xinput33 wbs_adr_i[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xinput44 wbs_dat_i[18] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_4
XFILLER_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput55 wbs_dat_i[28] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput66 wbs_dat_i[9] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
XFILLER_200_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1226_ net43 spm.x\[17\] _0410_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1157_ _0911_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1088_ _0875_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2060_ clknet_leaf_27_wb_clk_i _0347_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_2
XFILLER_94_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1011_ net40 Y\[14\] _0821_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__mux2_1
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ clknet_leaf_17_wb_clk_i _0002_ _0046_ VGND VGND VPWR VPWR spm.genblk1\[11\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1844_ _0592_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__buf_4
XFILLER_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1775_ _0614_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__clkbuf_4
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2327_ net143 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_111_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ net52 spm.x\[25\] _0399_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux2_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1560_ _0589_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
XFILLER_193_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1491_ _0583_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_193_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2112_ clknet_leaf_11_wb_clk_i spm.genblk1\[28\].csa.hsum2 _0212_ VGND VGND VPWR
+ VPWR spm.genblk1\[27\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ clknet_leaf_28_wb_clk_i _0330_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_2
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1827_ _0787_ _0749_ _0750_ _0606_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__a211o_1
XFILLER_117_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1758_ net115 _0657_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__and2_1
XFILLER_117_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1689_ P0\[37\] _0612_ _0615_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__o21a_1
XFILLER_85_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0991_ net47 Y\[20\] _0799_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__mux2_1
XFILLER_146_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1612_ _0595_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
XFILLER_114_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1543_ _0588_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1474_ _0574_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nor2_1
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2026_ clknet_leaf_27_wb_clk_i _0313_ _0159_ VGND VGND VPWR VPWR P0\[47\] sky130_fd_sc_hd__dfrtp_1
XFILLER_165_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1190_ _0928_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 wbs_adr_i[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0974_ _0802_ Y\[27\] _0794_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux2_1
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1526_ _0586_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1457_ _0452_ spm.x\[22\] VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1388_ spm.genblk1\[1\].csa.sc spm.genblk1\[1\].csa.y VGND VGND VPWR VPWR _0518_
+ sky130_fd_sc_hd__nor2_1
XSPM_example_150 VGND VGND VPWR VPWR SPM_example_150/HI io_out[5] sky130_fd_sc_hd__conb_1
XSPM_example_161 VGND VGND VPWR VPWR SPM_example_161/HI io_out[16] sky130_fd_sc_hd__conb_1
XSPM_example_172 VGND VGND VPWR VPWR SPM_example_172/HI io_out[27] sky130_fd_sc_hd__conb_1
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_183 VGND VGND VPWR VPWR SPM_example_183/HI irq[0] sky130_fd_sc_hd__conb_1
XFILLER_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_194 VGND VGND VPWR VPWR SPM_example_194/HI la_data_out[8] sky130_fd_sc_hd__conb_1
XFILLER_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ clknet_leaf_10_wb_clk_i _0296_ _0142_ VGND VGND VPWR VPWR P0\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1311_ _0453_ spm.x\[14\] VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nand2_1
XFILLER_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1242_ _0423_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1173_ P0\[8\] P0\[9\] _0914_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__mux2_1
XFILLER_64_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_14 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_25 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_47 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_58 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0957_ net58 Y\[30\] _0786_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__mux2_1
XFILLER_203_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput110 net110 VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput121 net121 VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput132 net132 VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_86_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_wb_clk_i clknet_2_0__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1509_ _0585_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__inv_2
XFILLER_142_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ _0760_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__inv_2
XFILLER_203_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 wbs_adr_i[19] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
X_1791_ P0\[55\] _0708_ _0709_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__o21a_1
Xinput23 wbs_adr_i[29] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput34 wbs_cyc_i VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput45 wbs_dat_i[19] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_4
Xinput56 wbs_dat_i[29] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput67 wbs_stb_i VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1225_ _0414_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1156_ P0\[16\] P0\[17\] _0903_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__mux2_1
XFILLER_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1087_ P0\[49\] P0\[50\] _0870_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__mux2_1
XFILLER_34_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1989_ clknet_leaf_22_wb_clk_i _0276_ _0122_ VGND VGND VPWR VPWR P0\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_140_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1010_ _0827_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1912_ clknet_leaf_17_wb_clk_i spm.genblk1\[11\].csa.hsum2 _0045_ VGND VGND VPWR
+ VPWR spm.genblk1\[10\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_176_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1843_ _0598_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__inv_2
XFILLER_129_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1774_ _0611_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__clkbuf_4
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ net141 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1208_ _0405_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1139_ P0\[24\] P0\[25\] _0892_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__mux2_1
XFILLER_26_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1490_ _0583_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_165_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2111_ clknet_leaf_13_wb_clk_i _0021_ _0211_ VGND VGND VPWR VPWR spm.genblk1\[29\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2042_ clknet_leaf_10_wb_clk_i _0329_ _0175_ VGND VGND VPWR VPWR P0\[63\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1826_ Y\[30\] _0778_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__and2_1
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1757_ P0\[49\] _0661_ _0662_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o21a_1
XFILLER_102_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1688_ Y\[5\] _0779_ _0635_ _0636_ _0606_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__a221o_1
XFILLER_172_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ net141 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_161_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0990_ _0813_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1611_ _0595_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__inv_2
XFILLER_154_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1542_ _0588_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
XFILLER_114_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1473_ spm.genblk1\[19\].csa.sc spm.genblk1\[19\].csa.y VGND VGND VPWR VPWR _0575_
+ sky130_fd_sc_hd__and2_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_310 VGND VGND VPWR VPWR SPM_example_310/HI la_data_out[124] sky130_fd_sc_hd__conb_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2025_ clknet_leaf_26_wb_clk_i _0312_ _0158_ VGND VGND VPWR VPWR P0\[46\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1809_ spm.x\[27\] P0\[27\] _0398_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__mux2_1
XFILLER_102_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0973_ net53 Y\[26\] _0799_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__mux2_1
XFILLER_146_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1525_ _0586_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__inv_2
XFILLER_82_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1456_ _0562_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__nor2_1
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1387_ _0497_ spm.x\[2\] _0516_ _0515_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__a31o_1
XSPM_example_151 VGND VGND VPWR VPWR SPM_example_151/HI io_out[6] sky130_fd_sc_hd__conb_1
XFILLER_68_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_162 VGND VGND VPWR VPWR SPM_example_162/HI io_out[17] sky130_fd_sc_hd__conb_1
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_173 VGND VGND VPWR VPWR SPM_example_173/HI io_out[28] sky130_fd_sc_hd__conb_1
XSPM_example_184 VGND VGND VPWR VPWR SPM_example_184/HI irq[1] sky130_fd_sc_hd__conb_1
XSPM_example_195 VGND VGND VPWR VPWR SPM_example_195/HI la_data_out[9] sky130_fd_sc_hd__conb_1
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2008_ clknet_leaf_9_wb_clk_i _0295_ _0141_ VGND VGND VPWR VPWR P0\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_211_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ _0464_ _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__nor2_1
XFILLER_123_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1241_ net36 spm.x\[10\] _0421_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1172_ _0919_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_37 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_59 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0956_ Y\[31\] _0779_ _0789_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o21a_1
XFILLER_146_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput100 net100 VGND VGND VPWR VPWR io_oeb[4] sky130_fd_sc_hd__buf_2
Xoutput111 net111 VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput122 net122 VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput133 net133 VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_47_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1508_ _0585_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__inv_2
XFILLER_102_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1439_ _0521_ spm.x\[25\] VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nand2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 wbs_adr_i[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_1790_ Y\[23\] _0700_ _0682_ _0720_ _0692_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__a221o_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput24 wbs_adr_i[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xinput35 wbs_dat_i[0] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_4
XFILLER_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput46 wbs_dat_i[1] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_4
Xinput57 wbs_dat_i[2] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput68 wbs_we_i VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
XFILLER_115_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1224_ net44 spm.x\[18\] _0410_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1155_ _0910_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1086_ _0874_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ clknet_leaf_22_wb_clk_i _0275_ _0121_ VGND VGND VPWR VPWR P0\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_165_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0939_ net15 net14 net17 net16 VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__or4_1
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ clknet_leaf_22_wb_clk_i _0003_ _0044_ VGND VGND VPWR VPWR spm.genblk1\[12\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_203_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1842_ _0598_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__inv_2
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1773_ Y\[20\] _0700_ _0682_ _0706_ _0692_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__a221o_1
XFILLER_184_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ net143 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1207_ net53 spm.x\[26\] _0399_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_1
XFILLER_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1138_ _0901_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1069_ _0865_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clknet_2_3__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_191_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2110_ clknet_leaf_13_wb_clk_i spm.genblk1\[29\].csa.hsum2 _0210_ VGND VGND VPWR
+ VPWR spm.genblk1\[28\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2041_ clknet_leaf_10_wb_clk_i _0328_ _0174_ VGND VGND VPWR VPWR P0\[62\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1825_ spm.x\[30\] P0\[30\] _0398_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__mux2_1
XFILLER_209_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1756_ Y\[17\] _0653_ _0682_ _0691_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__a221o_1
XFILLER_116_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1687_ spm.x\[5\] P0\[5\] _0622_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux2_1
XFILLER_116_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ net141 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1610_ _0595_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
XFILLER_201_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1541_ _0588_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
XFILLER_153_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1472_ spm.genblk1\[19\].csa.sc spm.genblk1\[19\].csa.y VGND VGND VPWR VPWR _0574_
+ sky130_fd_sc_hd__nor2_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_300 VGND VGND VPWR VPWR SPM_example_300/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_311 VGND VGND VPWR VPWR SPM_example_311/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XFILLER_39_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2024_ clknet_leaf_26_wb_clk_i _0311_ _0157_ VGND VGND VPWR VPWR P0\[45\] sky130_fd_sc_hd__dfrtp_1
XFILLER_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1808_ _0733_ _0734_ _0735_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a21o_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1739_ Y\[14\] _0653_ _0635_ _0678_ _0645_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__a221o_1
XFILLER_132_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0972_ _0801_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1524_ _0586_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__inv_2
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1455_ spm.genblk1\[22\].csa.sc spm.genblk1\[22\].csa.y VGND VGND VPWR VPWR _0563_
+ sky130_fd_sc_hd__and2_1
XFILLER_101_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1386_ _0516_ _0517_ VGND VGND VPWR VPWR spm.genblk1\[2\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_56_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSPM_example_152 VGND VGND VPWR VPWR SPM_example_152/HI io_out[7] sky130_fd_sc_hd__conb_1
XSPM_example_163 VGND VGND VPWR VPWR SPM_example_163/HI io_out[18] sky130_fd_sc_hd__conb_1
XFILLER_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_174 VGND VGND VPWR VPWR SPM_example_174/HI io_out[29] sky130_fd_sc_hd__conb_1
XSPM_example_185 VGND VGND VPWR VPWR SPM_example_185/HI irq[2] sky130_fd_sc_hd__conb_1
XSPM_example_196 VGND VGND VPWR VPWR SPM_example_196/HI la_data_out[10] sky130_fd_sc_hd__conb_1
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2007_ clknet_leaf_9_wb_clk_i _0294_ _0140_ VGND VGND VPWR VPWR P0\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1240_ _0422_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1171_ P0\[9\] P0\[10\] _0914_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__mux2_1
XFILLER_38_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_16 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_27 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_38 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_49 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0955_ net59 _0787_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__o21ba_1
XFILLER_203_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR io_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_115_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput112 net112 VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_86_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput123 net123 VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput134 net134 VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_115_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1507_ _0582_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__buf_4
XFILLER_47_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1438_ _0550_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__nor2_1
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1369_ _0497_ spm.x\[5\] _0504_ _0503_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a31o_1
XFILLER_110_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 wbs_adr_i[20] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
Xinput25 wbs_adr_i[30] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput36 wbs_dat_i[10] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
XFILLER_128_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput47 wbs_dat_i[20] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput58 wbs_dat_i[30] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
XFILLER_183_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1223_ _0413_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1154_ P0\[17\] P0\[18\] _0903_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__mux2_1
XFILLER_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1085_ P0\[50\] P0\[51\] _0870_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__mux2_1
XFILLER_80_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1987_ clknet_leaf_22_wb_clk_i _0274_ _0120_ VGND VGND VPWR VPWR P0\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0938_ _0769_ _0770_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__or3_1
XFILLER_180_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1910_ clknet_leaf_16_wb_clk_i spm.genblk1\[12\].csa.hsum2 _0043_ VGND VGND VPWR
+ VPWR spm.genblk1\[11\].csa.y sky130_fd_sc_hd__dfrtp_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1841_ _0598_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__inv_2
XFILLER_129_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1772_ spm.x\[20\] P0\[20\] _0669_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__mux2_1
XFILLER_129_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2324_ net139 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1206_ _0404_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1137_ P0\[25\] P0\[26\] _0892_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__mux2_1
XFILLER_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1068_ P0\[58\] P0\[59\] _0859_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2040_ clknet_leaf_9_wb_clk_i _0327_ _0173_ VGND VGND VPWR VPWR P0\[61\] sky130_fd_sc_hd__dfrtp_1
XFILLER_181_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1824_ _0746_ _0747_ _0748_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a21o_1
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1755_ _0605_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__buf_2
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1686_ _0786_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2307_ net143 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ _0582_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__buf_4
XFILLER_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1471_ _0541_ spm.x\[20\] _0572_ _0571_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a31o_1
XFILLER_114_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_301 VGND VGND VPWR VPWR SPM_example_301/HI la_data_out[115] sky130_fd_sc_hd__conb_1
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSPM_example_312 VGND VGND VPWR VPWR SPM_example_312/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2023_ clknet_leaf_26_wb_clk_i _0310_ _0156_ VGND VGND VPWR VPWR P0\[44\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1807_ net125 _0704_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__and2_1
XFILLER_163_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1738_ spm.x\[14\] P0\[14\] _0669_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__mux2_1
XFILLER_102_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1669_ _0619_ _0620_ _0621_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a21o_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0971_ _0800_ Y\[28\] _0794_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1523_ _0586_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__inv_2
XFILLER_153_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1454_ spm.genblk1\[22\].csa.sc spm.genblk1\[22\].csa.y VGND VGND VPWR VPWR _0562_
+ sky130_fd_sc_hd__nor2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1385_ _0479_ spm.x\[2\] VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__nand2_1
XFILLER_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSPM_example_153 VGND VGND VPWR VPWR SPM_example_153/HI io_out[8] sky130_fd_sc_hd__conb_1
XSPM_example_164 VGND VGND VPWR VPWR SPM_example_164/HI io_out[19] sky130_fd_sc_hd__conb_1
XFILLER_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_175 VGND VGND VPWR VPWR SPM_example_175/HI io_out[30] sky130_fd_sc_hd__conb_1
XFILLER_83_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_186 VGND VGND VPWR VPWR SPM_example_186/HI la_data_out[0] sky130_fd_sc_hd__conb_1
XSPM_example_197 VGND VGND VPWR VPWR SPM_example_197/HI la_data_out[11] sky130_fd_sc_hd__conb_1
XFILLER_167_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2006_ clknet_leaf_9_wb_clk_i _0293_ _0139_ VGND VGND VPWR VPWR P0\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1170_ _0918_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_17 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_39 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0954_ STATE VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__buf_2
XFILLER_146_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput102 net102 VGND VGND VPWR VPWR io_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput124 net124 VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_115_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput135 net135 VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_82_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1506_ _0584_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__inv_2
XFILLER_86_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1437_ spm.genblk1\[25\].csa.sc spm.genblk1\[25\].csa.y VGND VGND VPWR VPWR _0551_
+ sky130_fd_sc_hd__and2_1
X_1368_ _0504_ _0505_ VGND VGND VPWR VPWR spm.genblk1\[5\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1299_ _0453_ spm.x\[16\] VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__nand2_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput15 wbs_adr_i[21] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 wbs_adr_i[31] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_183_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput37 wbs_dat_i[11] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_4
Xinput48 wbs_dat_i[21] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
XFILLER_128_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput59 wbs_dat_i[31] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2340_ net141 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1222_ net45 spm.x\[19\] _0410_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
XFILLER_38_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1153_ _0909_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1084_ _0873_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ clknet_leaf_22_wb_clk_i _0273_ _0119_ VGND VGND VPWR VPWR P0\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_105_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0937_ net67 net34 VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__nand2_8
XFILLER_105_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1840_ _0598_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__inv_2
XFILLER_204_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1771_ _0702_ _0703_ _0705_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a21o_1
XFILLER_204_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2323_ net141 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1205_ net54 spm.x\[27\] _0399_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1136_ _0900_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1067_ _0864_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1969_ clknet_leaf_10_wb_clk_i _0265_ _0102_ VGND VGND VPWR VPWR spm.x\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_wb_clk_i clknet_2_2__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1823_ net128 _0602_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__and2_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1754_ spm.x\[17\] P0\[17\] _0669_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
XFILLER_129_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1685_ _0632_ _0633_ _0634_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__a21o_1
XFILLER_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ net143 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1119_ _0891_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2099_ clknet_leaf_6_wb_clk_i _0386_ _0199_ VGND VGND VPWR VPWR Y\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1470_ _0572_ _0573_ VGND VGND VPWR VPWR spm.genblk1\[20\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_45_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_302 VGND VGND VPWR VPWR SPM_example_302/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XFILLER_45_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_313 VGND VGND VPWR VPWR SPM_example_313/HI la_data_out[127] sky130_fd_sc_hd__conb_1
XFILLER_209_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2022_ clknet_leaf_26_wb_clk_i _0309_ _0155_ VGND VGND VPWR VPWR P0\[43\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1806_ P0\[58\] _0708_ _0709_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__o21a_1
XFILLER_163_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1737_ _0675_ _0676_ _0677_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a21o_1
XFILLER_85_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1668_ net118 _0603_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__and2_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1599_ _0594_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0970_ net54 Y\[27\] _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__mux2_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1522_ _0586_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__inv_2
XFILLER_114_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1453_ _0541_ spm.x\[23\] _0560_ _0559_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a31o_1
XFILLER_45_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1384_ _0514_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nor2_1
XFILLER_110_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_154 VGND VGND VPWR VPWR SPM_example_154/HI io_out[9] sky130_fd_sc_hd__conb_1
XSPM_example_165 VGND VGND VPWR VPWR SPM_example_165/HI io_out[20] sky130_fd_sc_hd__conb_1
XSPM_example_176 VGND VGND VPWR VPWR SPM_example_176/HI io_out[31] sky130_fd_sc_hd__conb_1
XFILLER_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_187 VGND VGND VPWR VPWR SPM_example_187/HI la_data_out[1] sky130_fd_sc_hd__conb_1
XFILLER_83_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_198 VGND VGND VPWR VPWR SPM_example_198/HI la_data_out[12] sky130_fd_sc_hd__conb_1
X_2005_ clknet_leaf_9_wb_clk_i _0292_ _0138_ VGND VGND VPWR VPWR P0\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_18 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_29 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0953_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__clkbuf_4
XFILLER_202_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR io_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput114 net114 VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput125 net125 VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput136 net136 VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_173_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1505_ _0584_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__inv_2
XFILLER_115_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1436_ spm.genblk1\[25\].csa.sc spm.genblk1\[25\].csa.y VGND VGND VPWR VPWR _0550_
+ sky130_fd_sc_hd__nor2_1
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1367_ _0479_ spm.x\[5\] VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__nand2_1
XFILLER_95_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1298_ _0456_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nor2_1
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_943 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 wbs_adr_i[22] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 wbs_adr_i[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 wbs_dat_i[12] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 wbs_dat_i[22] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
XFILLER_182_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1221_ _0412_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1152_ P0\[18\] P0\[19\] _0903_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__mux2_1
XFILLER_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1083_ P0\[51\] P0\[52\] _0870_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ clknet_leaf_22_wb_clk_i _0272_ _0118_ VGND VGND VPWR VPWR P0\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0936_ net29 net28 net31 net30 VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__or4_4
XFILLER_88_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1419_ _0537_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__nor2_1
XFILLER_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1770_ net117 _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__and2_1
XFILLER_200_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ net139 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1204_ _0403_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
X_1135_ P0\[26\] P0\[27\] _0892_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__mux2_1
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1066_ P0\[59\] P0\[60\] _0859_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1968_ clknet_leaf_10_wb_clk_i _0264_ _0101_ VGND VGND VPWR VPWR spm.x\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1899_ _0582_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__inv_2
XFILLER_147_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1822_ P0\[61\] _0708_ _0709_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__o21a_1
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1753_ _0688_ _0689_ _0690_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a21o_1
XFILLER_184_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1684_ net133 _0603_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__and2_1
XFILLER_131_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ net142 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1118_ P0\[34\] P0\[35\] _0881_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__mux2_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ clknet_leaf_5_wb_clk_i _0385_ _0198_ VGND VGND VPWR VPWR Y\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1049_ _0853_ Y\[3\] _0839_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__mux2_1
XFILLER_94_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_303 VGND VGND VPWR VPWR SPM_example_303/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2021_ clknet_leaf_24_wb_clk_i _0308_ _0154_ VGND VGND VPWR VPWR P0\[42\] sky130_fd_sc_hd__dfrtp_1
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1805_ Y\[26\] _0700_ _0786_ _0732_ _0692_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__a221o_1
XFILLER_129_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1736_ net111 _0657_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__and2_1
XFILLER_145_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1667_ P0\[33\] _0612_ _0615_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__o21a_1
XFILLER_116_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1598_ _0594_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
XFILLER_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1521_ _0586_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__inv_2
XFILLER_153_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1452_ _0560_ _0561_ VGND VGND VPWR VPWR spm.genblk1\[23\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1383_ spm.genblk1\[2\].csa.sc spm.genblk1\[2\].csa.y VGND VGND VPWR VPWR _0515_
+ sky130_fd_sc_hd__and2_1
XFILLER_171_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSPM_example_144 VGND VGND VPWR VPWR SPM_example_144/HI io_oeb[37] sky130_fd_sc_hd__conb_1
XFILLER_110_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSPM_example_155 VGND VGND VPWR VPWR SPM_example_155/HI io_out[10] sky130_fd_sc_hd__conb_1
XSPM_example_166 VGND VGND VPWR VPWR SPM_example_166/HI io_out[21] sky130_fd_sc_hd__conb_1
XFILLER_209_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_177 VGND VGND VPWR VPWR SPM_example_177/HI io_out[32] sky130_fd_sc_hd__conb_1
XSPM_example_188 VGND VGND VPWR VPWR SPM_example_188/HI la_data_out[2] sky130_fd_sc_hd__conb_1
XFILLER_55_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSPM_example_199 VGND VGND VPWR VPWR SPM_example_199/HI la_data_out[13] sky130_fd_sc_hd__conb_1
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2004_ clknet_leaf_7_wb_clk_i _0291_ _0137_ VGND VGND VPWR VPWR P0\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1719_ P0\[42\] _0661_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__o21a_1
XFILLER_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_19 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0952_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__clkbuf_4
XFILLER_159_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR io_oeb[8] sky130_fd_sc_hd__buf_2
Xoutput115 net115 VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_114_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput126 net126 VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput137 net137 VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__buf_2
X_1504_ _0584_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
XFILLER_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1435_ _0541_ spm.x\[26\] _0548_ _0547_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a31o_1
XFILLER_114_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1366_ _0502_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__nor2_1
XFILLER_56_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1297_ spm.genblk1\[16\].csa.sc spm.genblk1\[16\].csa.y VGND VGND VPWR VPWR _0457_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_15_wb_clk_i clknet_2_3__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 wbs_adr_i[23] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 wbs_adr_i[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
XFILLER_168_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput39 wbs_dat_i[13] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1220_ net47 spm.x\[20\] _0410_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1151_ _0908_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1082_ _0872_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1984_ clknet_leaf_21_wb_clk_i _0271_ _0117_ VGND VGND VPWR VPWR P0\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0935_ net68 VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__inv_2
XFILLER_14_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1418_ spm.genblk1\[28\].csa.sc spm.genblk1\[28\].csa.y VGND VGND VPWR VPWR _0538_
+ sky130_fd_sc_hd__and2_1
XFILLER_25_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1349_ _0491_ _0492_ VGND VGND VPWR VPWR spm.genblk1\[8\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1010 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ net139 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_152_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1203_ net55 spm.x\[28\] _0399_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux2_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1134_ _0899_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _0863_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1967_ clknet_leaf_11_wb_clk_i _0263_ _0100_ VGND VGND VPWR VPWR spm.x\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_105_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1898_ _0763_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__inv_2
XFILLER_107_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1821_ Y\[29\] _0700_ _0786_ _0745_ _0605_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a221o_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1752_ net114 _0657_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__and2_1
XFILLER_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1683_ P0\[36\] _0612_ _0615_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__o21a_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ net142 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1117_ _0890_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2097_ clknet_leaf_5_wb_clk_i _0384_ _0197_ VGND VGND VPWR VPWR Y\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_198_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1048_ net57 Y\[2\] _0798_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__mux2_1
XFILLER_80_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_972 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_304 VGND VGND VPWR VPWR SPM_example_304/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2020_ clknet_leaf_24_wb_clk_i _0307_ _0153_ VGND VGND VPWR VPWR P0\[41\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1804_ spm.x\[26\] P0\[26\] _0397_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__mux2_1
XFILLER_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1735_ P0\[45\] _0661_ _0662_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__o21a_1
XFILLER_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1666_ Y\[1\] _0779_ _0787_ _0618_ _0606_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__a221o_1
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1597_ _0594_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1520_ _0586_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__inv_2
XFILLER_142_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1451_ _0521_ spm.x\[23\] VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__nand2_1
XFILLER_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1382_ spm.genblk1\[2\].csa.sc spm.genblk1\[2\].csa.y VGND VGND VPWR VPWR _0514_
+ sky130_fd_sc_hd__nor2_1
XFILLER_45_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_145 VGND VGND VPWR VPWR SPM_example_145/HI io_out[0] sky130_fd_sc_hd__conb_1
XSPM_example_156 VGND VGND VPWR VPWR SPM_example_156/HI io_out[11] sky130_fd_sc_hd__conb_1
XSPM_example_167 VGND VGND VPWR VPWR SPM_example_167/HI io_out[22] sky130_fd_sc_hd__conb_1
XSPM_example_178 VGND VGND VPWR VPWR SPM_example_178/HI io_out[33] sky130_fd_sc_hd__conb_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_189 VGND VGND VPWR VPWR SPM_example_189/HI la_data_out[3] sky130_fd_sc_hd__conb_1
XFILLER_209_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2003_ clknet_leaf_7_wb_clk_i _0290_ _0136_ VGND VGND VPWR VPWR P0\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1718_ _0614_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__buf_2
XFILLER_145_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1649_ net106 _0603_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nor2_1
XFILLER_63_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0951_ _0764_ _0768_ _0772_ _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__or4_1
XFILLER_202_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput105 net105 VGND VGND VPWR VPWR io_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput116 net116 VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput127 net127 VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput138 net138 VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__buf_2
X_1503_ _0584_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XFILLER_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1434_ _0548_ _0549_ VGND VGND VPWR VPWR spm.genblk1\[26\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_96_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1365_ spm.genblk1\[5\].csa.sc spm.genblk1\[5\].csa.y VGND VGND VPWR VPWR _0503_
+ sky130_fd_sc_hd__and2_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1296_ spm.genblk1\[16\].csa.sc spm.genblk1\[16\].csa.y VGND VGND VPWR VPWR _0456_
+ sky130_fd_sc_hd__nor2_1
XFILLER_209_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 wbs_adr_i[24] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
XFILLER_210_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 wbs_adr_i[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1150_ P0\[19\] P0\[20\] _0903_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__mux2_1
XFILLER_93_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1081_ P0\[52\] P0\[53\] _0870_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__mux2_1
XFILLER_206_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1983_ clknet_leaf_20_wb_clk_i _0270_ _0116_ VGND VGND VPWR VPWR P0\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0934_ net27 _0765_ _0766_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__or4_1
XFILLER_53_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1417_ spm.genblk1\[28\].csa.sc spm.genblk1\[28\].csa.y VGND VGND VPWR VPWR _0537_
+ sky130_fd_sc_hd__nor2_1
XFILLER_130_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1348_ _0479_ spm.x\[8\] VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__nand2_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1279_ _0443_ _0444_ VGND VGND VPWR VPWR ncnt\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout140 net141 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_4
XFILLER_102_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ net142 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1202_ _0402_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1133_ P0\[27\] P0\[28\] _0892_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__mux2_1
XFILLER_38_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1064_ P0\[60\] P0\[61\] _0859_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__mux2_1
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clknet_2_0__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1966_ clknet_leaf_8_wb_clk_i _0262_ _0099_ VGND VGND VPWR VPWR spm.x\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_144_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1897_ _0763_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__inv_2
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1820_ spm.x\[29\] P0\[29\] _0397_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__mux2_1
XFILLER_54_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1751_ P0\[48\] _0661_ _0662_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__o21a_1
XFILLER_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1682_ Y\[4\] _0779_ _0787_ _0631_ _0606_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__a221o_1
XFILLER_209_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1116_ P0\[35\] P0\[36\] _0881_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__mux2_1
XFILLER_54_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2096_ clknet_leaf_5_wb_clk_i _0383_ _0196_ VGND VGND VPWR VPWR Y\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1047_ _0852_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1949_ clknet_leaf_22_wb_clk_i _0245_ _0082_ VGND VGND VPWR VPWR spm.x\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1007 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_305 VGND VGND VPWR VPWR SPM_example_305/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XFILLER_80_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1803_ _0729_ _0730_ _0731_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a21o_1
XFILLER_176_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1734_ Y\[13\] _0653_ _0635_ _0674_ _0645_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__a221o_1
XFILLER_129_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1665_ spm.x\[1\] P0\[1\] _0398_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__mux2_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1596_ _0592_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__buf_4
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2079_ clknet_leaf_21_wb_clk_i _0366_ _0179_ VGND VGND VPWR VPWR Y\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1450_ _0558_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__nor2_1
XFILLER_206_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1381_ _0497_ spm.x\[3\] _0512_ _0511_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__a31o_1
XFILLER_150_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_146 VGND VGND VPWR VPWR SPM_example_146/HI io_out[1] sky130_fd_sc_hd__conb_1
XFILLER_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_157 VGND VGND VPWR VPWR SPM_example_157/HI io_out[12] sky130_fd_sc_hd__conb_1
XSPM_example_168 VGND VGND VPWR VPWR SPM_example_168/HI io_out[23] sky130_fd_sc_hd__conb_1
XSPM_example_179 VGND VGND VPWR VPWR SPM_example_179/HI io_out[34] sky130_fd_sc_hd__conb_1
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2002_ clknet_leaf_3_wb_clk_i _0289_ _0135_ VGND VGND VPWR VPWR P0\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1717_ _0611_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__clkbuf_4
XFILLER_160_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1648_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1579_ _0591_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0950_ _0780_ _0781_ _0782_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__or4_1
XFILLER_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput106 net106 VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput117 net117 VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_127_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput128 net128 VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_1502_ _0584_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_2
XFILLER_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1433_ _0521_ spm.x\[26\] VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__nand2_1
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1364_ spm.genblk1\[5\].csa.sc spm.genblk1\[5\].csa.y VGND VGND VPWR VPWR _0502_
+ sky130_fd_sc_hd__nor2_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1295_ _0455_ spm.x\[17\] _0451_ _0450_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a31o_1
XFILLER_3_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clknet_2_0__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 wbs_adr_i[25] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_122_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1080_ _0871_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1982_ clknet_leaf_20_wb_clk_i _0269_ _0115_ VGND VGND VPWR VPWR P0\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0933_ net33 net32 net4 net3 VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__or4_1
XFILLER_174_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1416_ _0497_ spm.x\[29\] _0535_ _0534_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__a31o_1
XFILLER_60_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1347_ _0489_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__nor2_1
XFILLER_112_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1278_ CNT\[4\] _0441_ _0788_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__o21ai_1
XFILLER_3_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout141 net1 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_6
XFILLER_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1201_ net56 spm.x\[29\] _0399_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux2_1
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1132_ _0898_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1063_ _0862_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1965_ clknet_leaf_8_wb_clk_i _0261_ _0098_ VGND VGND VPWR VPWR spm.x\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_105_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1896_ _0763_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__inv_2
XFILLER_105_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1750_ Y\[16\] _0653_ _0682_ _0687_ _0645_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a221o_1
XFILLER_15_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1681_ spm.x\[4\] P0\[4\] _0622_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__mux2_1
XFILLER_128_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1115_ _0889_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2095_ clknet_leaf_3_wb_clk_i _0382_ _0195_ VGND VGND VPWR VPWR Y\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1046_ _0851_ Y\[4\] _0839_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__mux2_1
XFILLER_81_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1948_ clknet_leaf_17_wb_clk_i _0244_ _0081_ VGND VGND VPWR VPWR spm.x\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_162_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1879_ _0762_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__inv_2
XFILLER_162_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_306 VGND VGND VPWR VPWR SPM_example_306/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XFILLER_192_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1802_ net124 _0704_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__and2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1733_ spm.x\[13\] P0\[13\] _0669_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__mux2_1
XFILLER_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1664_ _0607_ _0616_ _0617_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__a21o_1
XFILLER_176_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1595_ _0593_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
XFILLER_113_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ clknet_leaf_20_wb_clk_i _0365_ _0178_ VGND VGND VPWR VPWR Y\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1029_ _0840_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380_ _0512_ _0513_ VGND VGND VPWR VPWR spm.genblk1\[3\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_171_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_147 VGND VGND VPWR VPWR SPM_example_147/HI io_out[2] sky130_fd_sc_hd__conb_1
XFILLER_110_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSPM_example_158 VGND VGND VPWR VPWR SPM_example_158/HI io_out[13] sky130_fd_sc_hd__conb_1
XSPM_example_169 VGND VGND VPWR VPWR SPM_example_169/HI io_out[24] sky130_fd_sc_hd__conb_1
XFILLER_208_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2001_ clknet_leaf_5_wb_clk_i _0288_ _0134_ VGND VGND VPWR VPWR P0\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1716_ Y\[10\] _0653_ _0635_ _0659_ _0645_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__a221o_1
XFILLER_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1647_ _0768_ _0772_ _0777_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__o31a_2
XFILLER_160_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1578_ _0591_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_154_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput107 net107 VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_126_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput118 net118 VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_142_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput129 net129 VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__buf_2
X_1501_ _0584_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_2
XFILLER_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1432_ _0546_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__nor2_1
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1363_ _0497_ spm.x\[6\] _0500_ _0499_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a31o_1
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1294_ _0453_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ clknet_leaf_20_wb_clk_i _0268_ _0114_ VGND VGND VPWR VPWR P0\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0932_ net13 net2 VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__or2_4
XFILLER_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1415_ _0535_ _0536_ VGND VGND VPWR VPWR spm.genblk1\[29\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1346_ spm.genblk1\[8\].csa.sc spm.genblk1\[8\].csa.y VGND VGND VPWR VPWR _0490_
+ sky130_fd_sc_hd__and2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1277_ CNT\[3\] CNT\[4\] _0438_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and3_1
XFILLER_37_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout142 net143 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_6
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1200_ _0401_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1131_ P0\[28\] P0\[29\] _0892_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__mux2_1
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1062_ P0\[61\] P0\[62\] _0859_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__mux2_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1964_ clknet_leaf_7_wb_clk_i _0260_ _0097_ VGND VGND VPWR VPWR spm.x\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1895_ _0763_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
XFILLER_88_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1329_ _0452_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_4
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1680_ _0628_ _0629_ _0630_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a21o_1
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1012 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_983 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1114_ P0\[36\] P0\[37\] _0881_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__mux2_1
XFILLER_4_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2094_ clknet_leaf_4_wb_clk_i _0381_ _0194_ VGND VGND VPWR VPWR Y\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1045_ net60 Y\[3\] _0798_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__mux2_1
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1947_ clknet_leaf_17_wb_clk_i _0243_ _0080_ VGND VGND VPWR VPWR spm.x\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_175_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1878_ _0762_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__inv_2
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSPM_example_307 VGND VGND VPWR VPWR SPM_example_307/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XFILLER_0_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1801_ P0\[57\] _0708_ _0709_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__o21a_1
XFILLER_157_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ _0671_ _0672_ _0673_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a21o_1
XFILLER_157_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1663_ net107 _0603_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__and2_1
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1594_ _0593_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2077_ clknet_leaf_16_wb_clk_i _0364_ _0177_ VGND VGND VPWR VPWR Y\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_121_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1028_ _0838_ Y\[10\] _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__mux2_1
XFILLER_210_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clknet_2_2__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_148 VGND VGND VPWR VPWR SPM_example_148/HI io_out[3] sky130_fd_sc_hd__conb_1
XSPM_example_159 VGND VGND VPWR VPWR SPM_example_159/HI io_out[14] sky130_fd_sc_hd__conb_1
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2000_ clknet_leaf_5_wb_clk_i _0287_ _0133_ VGND VGND VPWR VPWR P0\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1715_ spm.x\[10\] P0\[10\] _0622_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux2_1
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1646_ _0929_ _0777_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or3_1
XFILLER_160_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1577_ _0591_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
XFILLER_113_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2129_ clknet_leaf_11_wb_clk_i _0012_ _0229_ VGND VGND VPWR VPWR spm.genblk1\[20\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1500_ _0584_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_2
Xoutput108 net108 VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput119 net119 VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1431_ spm.genblk1\[26\].csa.sc spm.genblk1\[26\].csa.y VGND VGND VPWR VPWR _0547_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1362_ _0500_ _0501_ VGND VGND VPWR VPWR spm.genblk1\[6\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput90 net90 VGND VGND VPWR VPWR io_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1293_ _0451_ _0454_ VGND VGND VPWR VPWR spm.genblk1\[17\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1629_ _0592_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__buf_4
XFILLER_121_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ clknet_leaf_22_wb_clk_i _0267_ _0113_ VGND VGND VPWR VPWR P0\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0931_ net6 net5 net8 net7 VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__or4_2
XFILLER_144_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1414_ _0521_ spm.x\[29\] VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nand2_1
XFILLER_151_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1345_ spm.genblk1\[8\].csa.sc spm.genblk1\[8\].csa.y VGND VGND VPWR VPWR _0489_
+ sky130_fd_sc_hd__nor2_1
XFILLER_151_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1276_ _0441_ _0442_ VGND VGND VPWR VPWR ncnt\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_209_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout143 net1 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_8
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1130_ _0897_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1061_ _0861_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ clknet_leaf_7_wb_clk_i _0259_ _0096_ VGND VGND VPWR VPWR spm.x\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1894_ _0763_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__inv_2
XFILLER_179_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1328_ _0476_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__nor2_1
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1259_ net46 spm.x\[1\] _0398_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_72_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1113_ _0888_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2093_ clknet_leaf_4_wb_clk_i _0380_ _0193_ VGND VGND VPWR VPWR Y\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1044_ _0850_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1946_ clknet_leaf_17_wb_clk_i _0242_ _0079_ VGND VGND VPWR VPWR spm.x\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1877_ _0592_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__buf_4
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_308 VGND VGND VPWR VPWR SPM_example_308/HI la_data_out[122] sky130_fd_sc_hd__conb_1
XFILLER_48_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1800_ Y\[25\] _0700_ _0786_ _0728_ _0692_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__a221o_1
XFILLER_15_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1731_ net110 _0657_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__and2_1
XFILLER_89_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1662_ P0\[32\] _0612_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__o21a_1
XFILLER_176_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1593_ _0593_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
XFILLER_98_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2076_ clknet_leaf_16_wb_clk_i _0363_ _0176_ VGND VGND VPWR VPWR spm.y sky130_fd_sc_hd__dfrtp_1
XFILLER_208_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1027_ _0793_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1929_ clknet_leaf_19_wb_clk_i _0024_ _0062_ VGND VGND VPWR VPWR spm.genblk1\[3\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSPM_example_149 VGND VGND VPWR VPWR SPM_example_149/HI io_out[4] sky130_fd_sc_hd__conb_1
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1714_ _0655_ _0656_ _0658_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__a21o_1
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1645_ net68 _0599_ _0770_ _0771_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__or4_1
XFILLER_144_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1576_ _0591_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
XFILLER_116_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2128_ clknet_leaf_15_wb_clk_i spm.genblk1\[20\].csa.hsum2 _0228_ VGND VGND VPWR
+ VPWR spm.genblk1\[19\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_199_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2059_ clknet_leaf_27_wb_clk_i _0346_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_2
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_181_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1430_ spm.genblk1\[26\].csa.sc spm.genblk1\[26\].csa.y VGND VGND VPWR VPWR _0546_
+ sky130_fd_sc_hd__nor2_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1361_ _0479_ spm.x\[6\] VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__nand2_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput80 net80 VGND VGND VPWR VPWR io_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput91 net91 VGND VGND VPWR VPWR io_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_150_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1292_ _0453_ spm.x\[17\] VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__nand2_1
XFILLER_23_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1628_ _0596_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__inv_2
XFILLER_8_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1559_ _0589_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
XFILLER_143_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ net24 VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__inv_2
XFILLER_187_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1413_ _0533_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__nor2_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1344_ _0455_ spm.x\[9\] _0487_ _0486_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__a31o_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1275_ CNT\[3\] _0438_ _0788_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1060_ P0\[62\] P0\[63\] _0859_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_1
XFILLER_81_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ clknet_leaf_7_wb_clk_i _0258_ _0095_ VGND VGND VPWR VPWR spm.x\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_174_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1893_ _0763_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__inv_2
XFILLER_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1327_ spm.genblk1\[11\].csa.sc spm.genblk1\[11\].csa.y VGND VGND VPWR VPWR _0477_
+ sky130_fd_sc_hd__and2_1
XFILLER_112_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1258_ _0431_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1189_ P0\[0\] P0\[1\] _0793_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__mux2_1
XFILLER_80_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1112_ P0\[37\] P0\[38\] _0881_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__mux2_1
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2092_ clknet_leaf_0_wb_clk_i _0379_ _0192_ VGND VGND VPWR VPWR Y\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1043_ _0849_ Y\[5\] _0839_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1945_ clknet_leaf_18_wb_clk_i _0241_ _0078_ VGND VGND VPWR VPWR spm.x\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_119_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1876_ _0761_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__inv_2
XFILLER_174_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_309 VGND VGND VPWR VPWR SPM_example_309/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XFILLER_48_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1730_ P0\[44\] _0661_ _0662_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o21a_1
XFILLER_102_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1661_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__buf_2
XFILLER_176_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1592_ _0593_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
XFILLER_98_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2075_ clknet_leaf_10_wb_clk_i _0362_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_4
XFILLER_35_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1026_ net66 Y\[9\] _0821_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__mux2_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1928_ clknet_leaf_18_wb_clk_i spm.genblk1\[3\].csa.hsum2 _0061_ VGND VGND VPWR VPWR
+ spm.genblk1\[2\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_120_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1859_ _0760_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__inv_2
XFILLER_194_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clknet_2_0__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1713_ net138 _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__and2_1
XFILLER_118_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1644_ net27 VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__inv_2
XFILLER_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1575_ _0591_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
XFILLER_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2127_ clknet_leaf_11_wb_clk_i _0013_ _0227_ VGND VGND VPWR VPWR spm.genblk1\[21\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ clknet_leaf_26_wb_clk_i _0345_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_2
XFILLER_82_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1009_ _0826_ Y\[16\] _0817_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__mux2_1
XFILLER_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1360_ _0498_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__nor2_1
Xoutput70 net70 VGND VGND VPWR VPWR io_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput81 net81 VGND VGND VPWR VPWR io_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput92 net92 VGND VGND VPWR VPWR io_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_150_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1291_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__buf_2
XFILLER_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1627_ _0596_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__inv_2
XFILLER_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1558_ _0589_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
XFILLER_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1489_ _0583_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_80_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1412_ spm.genblk1\[29\].csa.sc spm.genblk1\[29\].csa.y VGND VGND VPWR VPWR _0534_
+ sky130_fd_sc_hd__and2_1
XFILLER_190_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1343_ _0487_ _0488_ VGND VGND VPWR VPWR spm.genblk1\[9\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1274_ CNT\[3\] _0438_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__and2_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0989_ _0812_ Y\[22\] _0794_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__mux2_1
XFILLER_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ clknet_leaf_7_wb_clk_i _0257_ _0094_ VGND VGND VPWR VPWR spm.x\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1892_ _0763_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__inv_2
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1326_ spm.genblk1\[11\].csa.sc spm.genblk1\[11\].csa.y VGND VGND VPWR VPWR _0476_
+ sky130_fd_sc_hd__nor2_1
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1257_ net57 spm.x\[2\] _0421_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1188_ _0927_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1111_ _0887_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2091_ clknet_leaf_0_wb_clk_i _0378_ _0191_ VGND VGND VPWR VPWR Y\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1042_ net61 Y\[4\] _0798_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__mux2_1
XFILLER_207_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1944_ clknet_leaf_19_wb_clk_i _0240_ _0077_ VGND VGND VPWR VPWR spm.x\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1875_ _0761_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__inv_2
XFILLER_119_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1309_ spm.genblk1\[14\].csa.sc spm.genblk1\[14\].csa.y VGND VGND VPWR VPWR _0465_
+ sky130_fd_sc_hd__and2_1
XFILLER_85_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1660_ net27 _0929_ _0613_ _0610_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__o31ai_4
XFILLER_176_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1591_ _0593_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
XFILLER_125_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2074_ clknet_leaf_9_wb_clk_i _0361_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_4
XFILLER_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1025_ _0837_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1927_ clknet_leaf_19_wb_clk_i _0025_ _0060_ VGND VGND VPWR VPWR spm.genblk1\[4\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1858_ _0760_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__inv_2
XFILLER_200_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1789_ spm.x\[23\] P0\[23\] _0397_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux2_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1712_ _0602_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__buf_2
XFILLER_117_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _0771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1643_ _0598_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__inv_2
XFILLER_133_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1574_ _0591_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
XFILLER_98_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2126_ clknet_leaf_11_wb_clk_i spm.genblk1\[21\].csa.hsum2 _0226_ VGND VGND VPWR
+ VPWR spm.genblk1\[20\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_187_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2057_ clknet_leaf_28_wb_clk_i _0344_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_4
XFILLER_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1008_ net41 Y\[15\] _0821_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__mux2_1
XFILLER_210_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput71 net71 VGND VGND VPWR VPWR io_oeb[11] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VGND VGND VPWR VPWR io_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VGND VGND VPWR VPWR io_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1290_ spm.y VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__buf_2
XFILLER_163_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1626_ _0596_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__inv_2
XFILLER_160_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1557_ _0589_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1488_ _0583_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
XFILLER_41_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2109_ clknet_leaf_15_wb_clk_i _0023_ _0209_ VGND VGND VPWR VPWR spm.genblk1\[30\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_wb_clk_i clknet_2_3__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1411_ spm.genblk1\[29\].csa.sc spm.genblk1\[29\].csa.y VGND VGND VPWR VPWR _0533_
+ sky130_fd_sc_hd__nor2_1
XFILLER_138_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1342_ _0479_ spm.x\[9\] VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__nand2_1
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1273_ _0440_ VGND VGND VPWR VPWR ncnt\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_111_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0988_ net48 Y\[21\] _0799_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__mux2_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1609_ _0595_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__inv_2
XFILLER_160_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSPM_example_290 VGND VGND VPWR VPWR SPM_example_290/HI la_data_out[104] sky130_fd_sc_hd__conb_1
XFILLER_167_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ clknet_leaf_7_wb_clk_i _0256_ _0093_ VGND VGND VPWR VPWR spm.x\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1891_ _0763_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__inv_2
XFILLER_147_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1325_ _0455_ spm.x\[12\] _0474_ _0473_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a31o_1
XFILLER_69_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1256_ _0430_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1187_ P0\[1\] P0\[2\] _0793_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__mux2_1
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ P0\[38\] P0\[39\] _0881_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__mux2_1
XFILLER_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2090_ clknet_leaf_0_wb_clk_i _0377_ _0190_ VGND VGND VPWR VPWR Y\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_171_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1041_ _0848_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1943_ clknet_leaf_20_wb_clk_i _0239_ _0076_ VGND VGND VPWR VPWR spm.x\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_148_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1874_ _0761_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__inv_2
XFILLER_174_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1308_ spm.genblk1\[14\].csa.sc spm.genblk1\[14\].csa.y VGND VGND VPWR VPWR _0464_
+ sky130_fd_sc_hd__nor2_1
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1239_ net37 spm.x\[11\] _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
XFILLER_77_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1590_ _0593_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
XFILLER_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2073_ clknet_leaf_9_wb_clk_i _0360_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_2
XFILLER_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1024_ _0836_ Y\[11\] _0817_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__mux2_1
XFILLER_207_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1926_ clknet_leaf_19_wb_clk_i spm.genblk1\[4\].csa.hsum2 _0059_ VGND VGND VPWR VPWR
+ spm.genblk1\[3\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1857_ _0760_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__inv_2
XFILLER_135_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1788_ _0717_ _0718_ _0719_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a21o_1
XFILLER_200_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1711_ P0\[41\] _0612_ _0615_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__o21a_1
XFILLER_172_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_2 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ _0598_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__inv_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1573_ _0582_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__buf_4
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2125_ clknet_leaf_12_wb_clk_i _0014_ _0225_ VGND VGND VPWR VPWR spm.genblk1\[22\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2056_ clknet_leaf_24_wb_clk_i _0343_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_4
XFILLER_70_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1007_ _0825_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1909_ clknet_leaf_23_wb_clk_i _0004_ _0042_ VGND VGND VPWR VPWR spm.genblk1\[13\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput72 net72 VGND VGND VPWR VPWR io_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput83 net83 VGND VGND VPWR VPWR io_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput94 net94 VGND VGND VPWR VPWR io_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1625_ _0596_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__inv_2
XFILLER_126_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1556_ _0589_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1487_ _0583_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
XFILLER_80_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ clknet_leaf_13_wb_clk_i spm.genblk1\[30\].csa.hsum2 _0208_ VGND VGND VPWR
+ VPWR spm.genblk1\[29\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2039_ clknet_leaf_5_wb_clk_i _0326_ _0172_ VGND VGND VPWR VPWR P0\[60\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410_ _0497_ spm.x\[30\] _0531_ _0530_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a31o_1
XFILLER_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1341_ _0485_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nor2_1
XFILLER_110_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1272_ _0438_ _0788_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__and3b_1
XFILLER_77_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0987_ _0811_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1608_ _0595_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__inv_2
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1539_ _0587_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
XFILLER_113_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSPM_example_280 VGND VGND VPWR VPWR SPM_example_280/HI la_data_out[94] sky130_fd_sc_hd__conb_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_291 VGND VGND VPWR VPWR SPM_example_291/HI la_data_out[105] sky130_fd_sc_hd__conb_1
XFILLER_167_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1890_ _0763_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__inv_2
XFILLER_186_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_922 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1324_ _0474_ _0475_ VGND VGND VPWR VPWR spm.genblk1\[12\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_97_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1255_ net60 spm.x\[3\] _0421_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
XFILLER_204_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1186_ _0926_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_947 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1040_ _0847_ Y\[6\] _0839_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__mux2_1
XFILLER_206_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1942_ clknet_leaf_20_wb_clk_i _0238_ _0075_ VGND VGND VPWR VPWR spm.x\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1873_ _0761_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__inv_2
XFILLER_31_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1307_ _0455_ spm.x\[15\] _0462_ _0461_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a31o_1
XFILLER_42_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1238_ _0398_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1169_ P0\[10\] P0\[11\] _0914_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2072_ clknet_leaf_4_wb_clk_i _0359_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_1
XFILLER_94_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1023_ net36 Y\[10\] _0821_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__mux2_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1925_ clknet_leaf_19_wb_clk_i _0026_ _0058_ VGND VGND VPWR VPWR spm.genblk1\[5\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_6_wb_clk_i clknet_2_1__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1856_ _0760_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__inv_2
XFILLER_190_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1787_ net121 _0704_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__and2_1
XFILLER_190_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2339_ net140 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1710_ Y\[9\] _0653_ _0635_ _0654_ _0645_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__a221o_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1641_ _0598_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__inv_2
XANTENNA_3 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1572_ _0590_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
XFILLER_67_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2124_ clknet_leaf_13_wb_clk_i spm.genblk1\[22\].csa.hsum2 _0224_ VGND VGND VPWR
+ VPWR spm.genblk1\[21\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2055_ clknet_leaf_26_wb_clk_i _0342_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_4
XFILLER_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ _0824_ Y\[17\] _0817_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__mux2_1
XFILLER_74_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1908_ clknet_leaf_23_wb_clk_i spm.genblk1\[13\].csa.hsum2 _0041_ VGND VGND VPWR
+ VPWR spm.genblk1\[12\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_124_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1839_ _0598_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__inv_2
XFILLER_194_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput73 net73 VGND VGND VPWR VPWR io_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_123_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput84 net84 VGND VGND VPWR VPWR io_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_95_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput95 net95 VGND VGND VPWR VPWR io_oeb[33] sky130_fd_sc_hd__buf_2
XFILLER_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1624_ _0596_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__inv_2
XFILLER_126_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1555_ _0589_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
XFILLER_125_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1486_ _0583_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_141_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2107_ clknet_leaf_10_wb_clk_i _0394_ _0207_ VGND VGND VPWR VPWR Y\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2038_ clknet_leaf_5_wb_clk_i _0325_ _0171_ VGND VGND VPWR VPWR P0\[59\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1340_ spm.genblk1\[9\].csa.sc spm.genblk1\[10\].csa.sum VGND VGND VPWR VPWR _0486_
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_20_wb_clk_i clknet_2_2__leaf_wb_clk_i VGND VGND VPWR VPWR clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1271_ CNT\[1\] CNT\[0\] CNT\[2\] VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__a21o_1
XFILLER_49_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0986_ _0810_ Y\[23\] _0794_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__mux2_1
XFILLER_118_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1607_ _0592_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__buf_4
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1538_ _0587_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_2
XFILLER_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1469_ _0452_ spm.x\[20\] VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__nand2_1
XFILLER_80_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_270 VGND VGND VPWR VPWR SPM_example_270/HI la_data_out[84] sky130_fd_sc_hd__conb_1
XFILLER_95_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSPM_example_281 VGND VGND VPWR VPWR SPM_example_281/HI la_data_out[95] sky130_fd_sc_hd__conb_1
XSPM_example_292 VGND VGND VPWR VPWR SPM_example_292/HI la_data_out[106] sky130_fd_sc_hd__conb_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1323_ _0453_ spm.x\[12\] VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__nand2_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1254_ _0429_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1185_ P0\[2\] P0\[3\] _0793_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__mux2_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0969_ _0798_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__buf_4
XFILLER_174_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1941_ clknet_leaf_20_wb_clk_i _0237_ _0074_ VGND VGND VPWR VPWR spm.x\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1872_ _0761_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__inv_2
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1306_ _0462_ _0463_ VGND VGND VPWR VPWR spm.genblk1\[15\].csa.hsum2 sky130_fd_sc_hd__xnor2_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1237_ _0420_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1168_ _0917_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1099_ _0793_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2071_ clknet_leaf_5_wb_clk_i _0358_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_4
XFILLER_94_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1022_ _0835_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1924_ clknet_leaf_19_wb_clk_i spm.genblk1\[5\].csa.hsum2 _0057_ VGND VGND VPWR VPWR
+ spm.genblk1\[4\].csa.y sky130_fd_sc_hd__dfrtp_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1855_ _0592_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__buf_4
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1786_ P0\[54\] _0708_ _0709_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__o21a_1
XFILLER_190_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2338_ net140 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1640_ _0592_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__clkbuf_8
XFILLER_177_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1571_ _0590_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2123_ clknet_leaf_11_wb_clk_i _0015_ _0223_ VGND VGND VPWR VPWR spm.genblk1\[23\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2054_ clknet_leaf_23_wb_clk_i _0341_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1005_ net42 Y\[16\] _0821_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__mux2_1
XFILLER_35_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1907_ clknet_leaf_23_wb_clk_i _0005_ _0040_ VGND VGND VPWR VPWR spm.genblk1\[14\].csa.sc
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1838_ _0598_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
XFILLER_190_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1769_ _0602_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__buf_2
XFILLER_190_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput74 net74 VGND VGND VPWR VPWR io_oeb[14] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VGND VGND VPWR VPWR io_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_123_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput96 net96 VGND VGND VPWR VPWR io_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1623_ _0596_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__inv_2
XFILLER_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1554_ _0589_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
XFILLER_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1485_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__buf_4
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
.ends

